version https://git-lfs.github.com/spec/v1
oid sha256:64f5182a5a2c93cdf1cd05b823ea4e2029b8cee8022940a7c6648bf05557dd21
size 165350
