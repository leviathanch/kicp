version https://git-lfs.github.com/spec/v1
oid sha256:3309152b6f787309fc5462ce191c8e76c71fd9e71c43f0e43ac6a64ac4494727
size 23161
