version https://git-lfs.github.com/spec/v1
oid sha256:78b57f0c93ca0ddc3caff5fc719244fd0851593d6b106a6eb5660e79d27126d2
size 23115
