magic
tech sky130A
magscale 1 2
timestamp 1685855751
<< obsli1 >>
rect 1104 2159 178848 177361
<< obsm1 >>
rect 934 892 179110 179308
<< metal2 >>
rect 2962 179200 3018 180000
rect 8574 179200 8630 180000
rect 14186 179200 14242 180000
rect 19798 179200 19854 180000
rect 25410 179200 25466 180000
rect 31022 179200 31078 180000
rect 36634 179200 36690 180000
rect 42246 179200 42302 180000
rect 47858 179200 47914 180000
rect 53470 179200 53526 180000
rect 59082 179200 59138 180000
rect 64694 179200 64750 180000
rect 70306 179200 70362 180000
rect 75918 179200 75974 180000
rect 81530 179200 81586 180000
rect 87142 179200 87198 180000
rect 92754 179200 92810 180000
rect 98366 179200 98422 180000
rect 103978 179200 104034 180000
rect 109590 179200 109646 180000
rect 115202 179200 115258 180000
rect 120814 179200 120870 180000
rect 126426 179200 126482 180000
rect 132038 179200 132094 180000
rect 137650 179200 137706 180000
rect 143262 179200 143318 180000
rect 148874 179200 148930 180000
rect 154486 179200 154542 180000
rect 160098 179200 160154 180000
rect 165710 179200 165766 180000
rect 171322 179200 171378 180000
rect 176934 179200 176990 180000
rect 12898 0 12954 800
rect 38566 0 38622 800
rect 64234 0 64290 800
rect 89902 0 89958 800
rect 115570 0 115626 800
rect 141238 0 141294 800
rect 166906 0 166962 800
<< obsm2 >>
rect 938 179144 2906 179330
rect 3074 179144 8518 179330
rect 8686 179144 14130 179330
rect 14298 179144 19742 179330
rect 19910 179144 25354 179330
rect 25522 179144 30966 179330
rect 31134 179144 36578 179330
rect 36746 179144 42190 179330
rect 42358 179144 47802 179330
rect 47970 179144 53414 179330
rect 53582 179144 59026 179330
rect 59194 179144 64638 179330
rect 64806 179144 70250 179330
rect 70418 179144 75862 179330
rect 76030 179144 81474 179330
rect 81642 179144 87086 179330
rect 87254 179144 92698 179330
rect 92866 179144 98310 179330
rect 98478 179144 103922 179330
rect 104090 179144 109534 179330
rect 109702 179144 115146 179330
rect 115314 179144 120758 179330
rect 120926 179144 126370 179330
rect 126538 179144 131982 179330
rect 132150 179144 137594 179330
rect 137762 179144 143206 179330
rect 143374 179144 148818 179330
rect 148986 179144 154430 179330
rect 154598 179144 160042 179330
rect 160210 179144 165654 179330
rect 165822 179144 171266 179330
rect 171434 179144 176878 179330
rect 177046 179144 179106 179330
rect 938 856 179106 179144
rect 938 800 12842 856
rect 13010 800 38510 856
rect 38678 800 64178 856
rect 64346 800 89846 856
rect 90014 800 115514 856
rect 115682 800 141182 856
rect 141350 800 166850 856
rect 167018 800 179106 856
<< metal3 >>
rect 0 176264 800 176384
rect 179200 176264 180000 176384
rect 0 170688 800 170808
rect 179200 170688 180000 170808
rect 0 165112 800 165232
rect 179200 165112 180000 165232
rect 0 159536 800 159656
rect 179200 159536 180000 159656
rect 0 153960 800 154080
rect 179200 153960 180000 154080
rect 0 148384 800 148504
rect 179200 148384 180000 148504
rect 0 142808 800 142928
rect 179200 142808 180000 142928
rect 0 137232 800 137352
rect 179200 137232 180000 137352
rect 0 131656 800 131776
rect 179200 131656 180000 131776
rect 0 126080 800 126200
rect 179200 126080 180000 126200
rect 0 120504 800 120624
rect 179200 120504 180000 120624
rect 0 114928 800 115048
rect 179200 114928 180000 115048
rect 0 109352 800 109472
rect 179200 109352 180000 109472
rect 0 103776 800 103896
rect 179200 103776 180000 103896
rect 0 98200 800 98320
rect 179200 98200 180000 98320
rect 0 92624 800 92744
rect 179200 92624 180000 92744
rect 0 87048 800 87168
rect 179200 87048 180000 87168
rect 0 81472 800 81592
rect 179200 81472 180000 81592
rect 0 75896 800 76016
rect 179200 75896 180000 76016
rect 0 70320 800 70440
rect 179200 70320 180000 70440
rect 0 64744 800 64864
rect 179200 64744 180000 64864
rect 0 59168 800 59288
rect 179200 59168 180000 59288
rect 0 53592 800 53712
rect 179200 53592 180000 53712
rect 0 48016 800 48136
rect 179200 48016 180000 48136
rect 0 42440 800 42560
rect 179200 42440 180000 42560
rect 0 36864 800 36984
rect 179200 36864 180000 36984
rect 0 31288 800 31408
rect 179200 31288 180000 31408
rect 0 25712 800 25832
rect 179200 25712 180000 25832
rect 0 20136 800 20256
rect 179200 20136 180000 20256
rect 0 14560 800 14680
rect 179200 14560 180000 14680
rect 0 8984 800 9104
rect 179200 8984 180000 9104
rect 0 3408 800 3528
rect 179200 3408 180000 3528
<< obsm3 >>
rect 800 176464 179200 177377
rect 880 176184 179120 176464
rect 800 170888 179200 176184
rect 880 170608 179120 170888
rect 800 165312 179200 170608
rect 880 165032 179120 165312
rect 800 159736 179200 165032
rect 880 159456 179120 159736
rect 800 154160 179200 159456
rect 880 153880 179120 154160
rect 800 148584 179200 153880
rect 880 148304 179120 148584
rect 800 143008 179200 148304
rect 880 142728 179120 143008
rect 800 137432 179200 142728
rect 880 137152 179120 137432
rect 800 131856 179200 137152
rect 880 131576 179120 131856
rect 800 126280 179200 131576
rect 880 126000 179120 126280
rect 800 120704 179200 126000
rect 880 120424 179120 120704
rect 800 115128 179200 120424
rect 880 114848 179120 115128
rect 800 109552 179200 114848
rect 880 109272 179120 109552
rect 800 103976 179200 109272
rect 880 103696 179120 103976
rect 800 98400 179200 103696
rect 880 98120 179120 98400
rect 800 92824 179200 98120
rect 880 92544 179120 92824
rect 800 87248 179200 92544
rect 880 86968 179120 87248
rect 800 81672 179200 86968
rect 880 81392 179120 81672
rect 800 76096 179200 81392
rect 880 75816 179120 76096
rect 800 70520 179200 75816
rect 880 70240 179120 70520
rect 800 64944 179200 70240
rect 880 64664 179120 64944
rect 800 59368 179200 64664
rect 880 59088 179120 59368
rect 800 53792 179200 59088
rect 880 53512 179120 53792
rect 800 48216 179200 53512
rect 880 47936 179120 48216
rect 800 42640 179200 47936
rect 880 42360 179120 42640
rect 800 37064 179200 42360
rect 880 36784 179120 37064
rect 800 31488 179200 36784
rect 880 31208 179120 31488
rect 800 25912 179200 31208
rect 880 25632 179120 25912
rect 800 20336 179200 25632
rect 880 20056 179120 20336
rect 800 14760 179200 20056
rect 880 14480 179120 14760
rect 800 9184 179200 14480
rect 880 8904 179120 9184
rect 800 3608 179200 8904
rect 880 3328 179120 3608
rect 800 2143 179200 3328
<< metal4 >>
rect 4208 2128 4528 177392
rect 19568 2128 19888 177392
rect 34928 2128 35248 177392
rect 50288 2128 50608 177392
rect 65648 2128 65968 177392
rect 81008 2128 81328 177392
rect 96368 2128 96688 177392
rect 111728 2128 112048 177392
rect 127088 2128 127408 177392
rect 142448 2128 142768 177392
rect 157808 2128 158128 177392
rect 173168 2128 173488 177392
<< obsm4 >>
rect 4659 2347 19488 176765
rect 19968 2347 34848 176765
rect 35328 2347 50208 176765
rect 50688 2347 65568 176765
rect 66048 2347 80928 176765
rect 81408 2347 96288 176765
rect 96768 2347 111648 176765
rect 112128 2347 127008 176765
rect 127488 2347 142368 176765
rect 142848 2347 157728 176765
rect 158208 2347 173088 176765
rect 173568 2347 174189 176765
<< labels >>
rlabel metal2 s 2962 179200 3018 180000 6 addr_o[0]
port 1 nsew signal output
rlabel metal2 s 59082 179200 59138 180000 6 addr_o[10]
port 2 nsew signal output
rlabel metal2 s 64694 179200 64750 180000 6 addr_o[11]
port 3 nsew signal output
rlabel metal2 s 70306 179200 70362 180000 6 addr_o[12]
port 4 nsew signal output
rlabel metal2 s 75918 179200 75974 180000 6 addr_o[13]
port 5 nsew signal output
rlabel metal2 s 81530 179200 81586 180000 6 addr_o[14]
port 6 nsew signal output
rlabel metal2 s 87142 179200 87198 180000 6 addr_o[15]
port 7 nsew signal output
rlabel metal2 s 92754 179200 92810 180000 6 addr_o[16]
port 8 nsew signal output
rlabel metal2 s 98366 179200 98422 180000 6 addr_o[17]
port 9 nsew signal output
rlabel metal2 s 103978 179200 104034 180000 6 addr_o[18]
port 10 nsew signal output
rlabel metal2 s 109590 179200 109646 180000 6 addr_o[19]
port 11 nsew signal output
rlabel metal2 s 8574 179200 8630 180000 6 addr_o[1]
port 12 nsew signal output
rlabel metal2 s 115202 179200 115258 180000 6 addr_o[20]
port 13 nsew signal output
rlabel metal2 s 120814 179200 120870 180000 6 addr_o[21]
port 14 nsew signal output
rlabel metal2 s 126426 179200 126482 180000 6 addr_o[22]
port 15 nsew signal output
rlabel metal2 s 132038 179200 132094 180000 6 addr_o[23]
port 16 nsew signal output
rlabel metal2 s 137650 179200 137706 180000 6 addr_o[24]
port 17 nsew signal output
rlabel metal2 s 143262 179200 143318 180000 6 addr_o[25]
port 18 nsew signal output
rlabel metal2 s 148874 179200 148930 180000 6 addr_o[26]
port 19 nsew signal output
rlabel metal2 s 154486 179200 154542 180000 6 addr_o[27]
port 20 nsew signal output
rlabel metal2 s 160098 179200 160154 180000 6 addr_o[28]
port 21 nsew signal output
rlabel metal2 s 165710 179200 165766 180000 6 addr_o[29]
port 22 nsew signal output
rlabel metal2 s 14186 179200 14242 180000 6 addr_o[2]
port 23 nsew signal output
rlabel metal2 s 171322 179200 171378 180000 6 addr_o[30]
port 24 nsew signal output
rlabel metal2 s 176934 179200 176990 180000 6 addr_o[31]
port 25 nsew signal output
rlabel metal2 s 19798 179200 19854 180000 6 addr_o[3]
port 26 nsew signal output
rlabel metal2 s 25410 179200 25466 180000 6 addr_o[4]
port 27 nsew signal output
rlabel metal2 s 31022 179200 31078 180000 6 addr_o[5]
port 28 nsew signal output
rlabel metal2 s 36634 179200 36690 180000 6 addr_o[6]
port 29 nsew signal output
rlabel metal2 s 42246 179200 42302 180000 6 addr_o[7]
port 30 nsew signal output
rlabel metal2 s 47858 179200 47914 180000 6 addr_o[8]
port 31 nsew signal output
rlabel metal2 s 53470 179200 53526 180000 6 addr_o[9]
port 32 nsew signal output
rlabel metal2 s 12898 0 12954 800 6 clk
port 33 nsew signal input
rlabel metal3 s 179200 3408 180000 3528 6 data_i[0]
port 34 nsew signal input
rlabel metal3 s 179200 59168 180000 59288 6 data_i[10]
port 35 nsew signal input
rlabel metal3 s 179200 64744 180000 64864 6 data_i[11]
port 36 nsew signal input
rlabel metal3 s 179200 70320 180000 70440 6 data_i[12]
port 37 nsew signal input
rlabel metal3 s 179200 75896 180000 76016 6 data_i[13]
port 38 nsew signal input
rlabel metal3 s 179200 81472 180000 81592 6 data_i[14]
port 39 nsew signal input
rlabel metal3 s 179200 87048 180000 87168 6 data_i[15]
port 40 nsew signal input
rlabel metal3 s 179200 92624 180000 92744 6 data_i[16]
port 41 nsew signal input
rlabel metal3 s 179200 98200 180000 98320 6 data_i[17]
port 42 nsew signal input
rlabel metal3 s 179200 103776 180000 103896 6 data_i[18]
port 43 nsew signal input
rlabel metal3 s 179200 109352 180000 109472 6 data_i[19]
port 44 nsew signal input
rlabel metal3 s 179200 8984 180000 9104 6 data_i[1]
port 45 nsew signal input
rlabel metal3 s 179200 114928 180000 115048 6 data_i[20]
port 46 nsew signal input
rlabel metal3 s 179200 120504 180000 120624 6 data_i[21]
port 47 nsew signal input
rlabel metal3 s 179200 126080 180000 126200 6 data_i[22]
port 48 nsew signal input
rlabel metal3 s 179200 131656 180000 131776 6 data_i[23]
port 49 nsew signal input
rlabel metal3 s 179200 137232 180000 137352 6 data_i[24]
port 50 nsew signal input
rlabel metal3 s 179200 142808 180000 142928 6 data_i[25]
port 51 nsew signal input
rlabel metal3 s 179200 148384 180000 148504 6 data_i[26]
port 52 nsew signal input
rlabel metal3 s 179200 153960 180000 154080 6 data_i[27]
port 53 nsew signal input
rlabel metal3 s 179200 159536 180000 159656 6 data_i[28]
port 54 nsew signal input
rlabel metal3 s 179200 165112 180000 165232 6 data_i[29]
port 55 nsew signal input
rlabel metal3 s 179200 14560 180000 14680 6 data_i[2]
port 56 nsew signal input
rlabel metal3 s 179200 170688 180000 170808 6 data_i[30]
port 57 nsew signal input
rlabel metal3 s 179200 176264 180000 176384 6 data_i[31]
port 58 nsew signal input
rlabel metal3 s 179200 20136 180000 20256 6 data_i[3]
port 59 nsew signal input
rlabel metal3 s 179200 25712 180000 25832 6 data_i[4]
port 60 nsew signal input
rlabel metal3 s 179200 31288 180000 31408 6 data_i[5]
port 61 nsew signal input
rlabel metal3 s 179200 36864 180000 36984 6 data_i[6]
port 62 nsew signal input
rlabel metal3 s 179200 42440 180000 42560 6 data_i[7]
port 63 nsew signal input
rlabel metal3 s 179200 48016 180000 48136 6 data_i[8]
port 64 nsew signal input
rlabel metal3 s 179200 53592 180000 53712 6 data_i[9]
port 65 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 data_o[0]
port 66 nsew signal output
rlabel metal3 s 0 59168 800 59288 6 data_o[10]
port 67 nsew signal output
rlabel metal3 s 0 64744 800 64864 6 data_o[11]
port 68 nsew signal output
rlabel metal3 s 0 70320 800 70440 6 data_o[12]
port 69 nsew signal output
rlabel metal3 s 0 75896 800 76016 6 data_o[13]
port 70 nsew signal output
rlabel metal3 s 0 81472 800 81592 6 data_o[14]
port 71 nsew signal output
rlabel metal3 s 0 87048 800 87168 6 data_o[15]
port 72 nsew signal output
rlabel metal3 s 0 92624 800 92744 6 data_o[16]
port 73 nsew signal output
rlabel metal3 s 0 98200 800 98320 6 data_o[17]
port 74 nsew signal output
rlabel metal3 s 0 103776 800 103896 6 data_o[18]
port 75 nsew signal output
rlabel metal3 s 0 109352 800 109472 6 data_o[19]
port 76 nsew signal output
rlabel metal3 s 0 8984 800 9104 6 data_o[1]
port 77 nsew signal output
rlabel metal3 s 0 114928 800 115048 6 data_o[20]
port 78 nsew signal output
rlabel metal3 s 0 120504 800 120624 6 data_o[21]
port 79 nsew signal output
rlabel metal3 s 0 126080 800 126200 6 data_o[22]
port 80 nsew signal output
rlabel metal3 s 0 131656 800 131776 6 data_o[23]
port 81 nsew signal output
rlabel metal3 s 0 137232 800 137352 6 data_o[24]
port 82 nsew signal output
rlabel metal3 s 0 142808 800 142928 6 data_o[25]
port 83 nsew signal output
rlabel metal3 s 0 148384 800 148504 6 data_o[26]
port 84 nsew signal output
rlabel metal3 s 0 153960 800 154080 6 data_o[27]
port 85 nsew signal output
rlabel metal3 s 0 159536 800 159656 6 data_o[28]
port 86 nsew signal output
rlabel metal3 s 0 165112 800 165232 6 data_o[29]
port 87 nsew signal output
rlabel metal3 s 0 14560 800 14680 6 data_o[2]
port 88 nsew signal output
rlabel metal3 s 0 170688 800 170808 6 data_o[30]
port 89 nsew signal output
rlabel metal3 s 0 176264 800 176384 6 data_o[31]
port 90 nsew signal output
rlabel metal3 s 0 20136 800 20256 6 data_o[3]
port 91 nsew signal output
rlabel metal3 s 0 25712 800 25832 6 data_o[4]
port 92 nsew signal output
rlabel metal3 s 0 31288 800 31408 6 data_o[5]
port 93 nsew signal output
rlabel metal3 s 0 36864 800 36984 6 data_o[6]
port 94 nsew signal output
rlabel metal3 s 0 42440 800 42560 6 data_o[7]
port 95 nsew signal output
rlabel metal3 s 0 48016 800 48136 6 data_o[8]
port 96 nsew signal output
rlabel metal3 s 0 53592 800 53712 6 data_o[9]
port 97 nsew signal output
rlabel metal2 s 115570 0 115626 800 6 done
port 98 nsew signal output
rlabel metal2 s 64234 0 64290 800 6 enable
port 99 nsew signal input
rlabel metal2 s 89902 0 89958 800 6 mem_opdone
port 100 nsew signal input
rlabel metal2 s 141238 0 141294 800 6 mem_operation[0]
port 101 nsew signal output
rlabel metal2 s 166906 0 166962 800 6 mem_operation[1]
port 102 nsew signal output
rlabel metal2 s 38566 0 38622 800 6 reset
port 103 nsew signal input
rlabel metal4 s 4208 2128 4528 177392 6 vccd1
port 104 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 177392 6 vccd1
port 104 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 177392 6 vccd1
port 104 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 177392 6 vccd1
port 104 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 177392 6 vccd1
port 104 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 177392 6 vccd1
port 104 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 177392 6 vssd1
port 105 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 177392 6 vssd1
port 105 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 177392 6 vssd1
port 105 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 177392 6 vssd1
port 105 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 177392 6 vssd1
port 105 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 177392 6 vssd1
port 105 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 180000 180000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 59634302
string GDS_FILE /home/leviathan/kicp/openlane/Matrix_Convolution/runs/23_06_04_05_03/results/signoff/Matrix_Convolution.magic.gds
string GDS_START 1526526
<< end >>

