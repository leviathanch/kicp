version https://git-lfs.github.com/spec/v1
oid sha256:33445ab1e2061708c7c87b5b001b8401023f5b4c5202cd77c448f6b7ac3d87c2
size 117602
