version https://git-lfs.github.com/spec/v1
oid sha256:b71ac77de1a3cc5c28fc23690b2631e7aeb66e3d5f02a209748f8069b9f05edf
size 23108
