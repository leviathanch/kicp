version https://git-lfs.github.com/spec/v1
oid sha256:4f9a941cbcdae748dd84b9901f118dda3858a3890d057592a39747033eb338d6
size 116385
