VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Matrix_Multiplication
  CLASS BLOCK ;
  FOREIGN Matrix_Multiplication ;
  ORIGIN 0.000 0.000 ;
  SIZE 900.000 BY 900.000 ;
  PIN addr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.810 896.000 15.090 900.000 ;
    END
  END addr_o[0]
  PIN addr_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.410 896.000 295.690 900.000 ;
    END
  END addr_o[10]
  PIN addr_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.470 896.000 323.750 900.000 ;
    END
  END addr_o[11]
  PIN addr_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.530 896.000 351.810 900.000 ;
    END
  END addr_o[12]
  PIN addr_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.590 896.000 379.870 900.000 ;
    END
  END addr_o[13]
  PIN addr_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.650 896.000 407.930 900.000 ;
    END
  END addr_o[14]
  PIN addr_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 435.710 896.000 435.990 900.000 ;
    END
  END addr_o[15]
  PIN addr_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.770 896.000 464.050 900.000 ;
    END
  END addr_o[16]
  PIN addr_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.830 896.000 492.110 900.000 ;
    END
  END addr_o[17]
  PIN addr_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.890 896.000 520.170 900.000 ;
    END
  END addr_o[18]
  PIN addr_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.950 896.000 548.230 900.000 ;
    END
  END addr_o[19]
  PIN addr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 896.000 43.150 900.000 ;
    END
  END addr_o[1]
  PIN addr_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.010 896.000 576.290 900.000 ;
    END
  END addr_o[20]
  PIN addr_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.070 896.000 604.350 900.000 ;
    END
  END addr_o[21]
  PIN addr_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.130 896.000 632.410 900.000 ;
    END
  END addr_o[22]
  PIN addr_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.190 896.000 660.470 900.000 ;
    END
  END addr_o[23]
  PIN addr_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.250 896.000 688.530 900.000 ;
    END
  END addr_o[24]
  PIN addr_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 716.310 896.000 716.590 900.000 ;
    END
  END addr_o[25]
  PIN addr_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 744.370 896.000 744.650 900.000 ;
    END
  END addr_o[26]
  PIN addr_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 772.430 896.000 772.710 900.000 ;
    END
  END addr_o[27]
  PIN addr_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.490 896.000 800.770 900.000 ;
    END
  END addr_o[28]
  PIN addr_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 828.550 896.000 828.830 900.000 ;
    END
  END addr_o[29]
  PIN addr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 896.000 71.210 900.000 ;
    END
  END addr_o[2]
  PIN addr_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 856.610 896.000 856.890 900.000 ;
    END
  END addr_o[30]
  PIN addr_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 884.670 896.000 884.950 900.000 ;
    END
  END addr_o[31]
  PIN addr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.990 896.000 99.270 900.000 ;
    END
  END addr_o[3]
  PIN addr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.050 896.000 127.330 900.000 ;
    END
  END addr_o[4]
  PIN addr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.110 896.000 155.390 900.000 ;
    END
  END addr_o[5]
  PIN addr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.170 896.000 183.450 900.000 ;
    END
  END addr_o[6]
  PIN addr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.230 896.000 211.510 900.000 ;
    END
  END addr_o[7]
  PIN addr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.290 896.000 239.570 900.000 ;
    END
  END addr_o[8]
  PIN addr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 896.000 267.630 900.000 ;
    END
  END addr_o[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END clk
  PIN data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 17.040 900.000 17.640 ;
    END
  END data_i[0]
  PIN data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 295.840 900.000 296.440 ;
    END
  END data_i[10]
  PIN data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 323.720 900.000 324.320 ;
    END
  END data_i[11]
  PIN data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 351.600 900.000 352.200 ;
    END
  END data_i[12]
  PIN data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 379.480 900.000 380.080 ;
    END
  END data_i[13]
  PIN data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 407.360 900.000 407.960 ;
    END
  END data_i[14]
  PIN data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 435.240 900.000 435.840 ;
    END
  END data_i[15]
  PIN data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 463.120 900.000 463.720 ;
    END
  END data_i[16]
  PIN data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 491.000 900.000 491.600 ;
    END
  END data_i[17]
  PIN data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 518.880 900.000 519.480 ;
    END
  END data_i[18]
  PIN data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 546.760 900.000 547.360 ;
    END
  END data_i[19]
  PIN data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 44.920 900.000 45.520 ;
    END
  END data_i[1]
  PIN data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 574.640 900.000 575.240 ;
    END
  END data_i[20]
  PIN data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 602.520 900.000 603.120 ;
    END
  END data_i[21]
  PIN data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 630.400 900.000 631.000 ;
    END
  END data_i[22]
  PIN data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 658.280 900.000 658.880 ;
    END
  END data_i[23]
  PIN data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 686.160 900.000 686.760 ;
    END
  END data_i[24]
  PIN data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 714.040 900.000 714.640 ;
    END
  END data_i[25]
  PIN data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 741.920 900.000 742.520 ;
    END
  END data_i[26]
  PIN data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 769.800 900.000 770.400 ;
    END
  END data_i[27]
  PIN data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 797.680 900.000 798.280 ;
    END
  END data_i[28]
  PIN data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 825.560 900.000 826.160 ;
    END
  END data_i[29]
  PIN data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 72.800 900.000 73.400 ;
    END
  END data_i[2]
  PIN data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 853.440 900.000 854.040 ;
    END
  END data_i[30]
  PIN data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 881.320 900.000 881.920 ;
    END
  END data_i[31]
  PIN data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 100.680 900.000 101.280 ;
    END
  END data_i[3]
  PIN data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 128.560 900.000 129.160 ;
    END
  END data_i[4]
  PIN data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 156.440 900.000 157.040 ;
    END
  END data_i[5]
  PIN data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 184.320 900.000 184.920 ;
    END
  END data_i[6]
  PIN data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 212.200 900.000 212.800 ;
    END
  END data_i[7]
  PIN data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 240.080 900.000 240.680 ;
    END
  END data_i[8]
  PIN data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 267.960 900.000 268.560 ;
    END
  END data_i[9]
  PIN data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END data_o[0]
  PIN data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.840 4.000 296.440 ;
    END
  END data_o[10]
  PIN data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.720 4.000 324.320 ;
    END
  END data_o[11]
  PIN data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 351.600 4.000 352.200 ;
    END
  END data_o[12]
  PIN data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 379.480 4.000 380.080 ;
    END
  END data_o[13]
  PIN data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 407.360 4.000 407.960 ;
    END
  END data_o[14]
  PIN data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.240 4.000 435.840 ;
    END
  END data_o[15]
  PIN data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 463.120 4.000 463.720 ;
    END
  END data_o[16]
  PIN data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 491.000 4.000 491.600 ;
    END
  END data_o[17]
  PIN data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 518.880 4.000 519.480 ;
    END
  END data_o[18]
  PIN data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 546.760 4.000 547.360 ;
    END
  END data_o[19]
  PIN data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 4.000 45.520 ;
    END
  END data_o[1]
  PIN data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 574.640 4.000 575.240 ;
    END
  END data_o[20]
  PIN data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 602.520 4.000 603.120 ;
    END
  END data_o[21]
  PIN data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 630.400 4.000 631.000 ;
    END
  END data_o[22]
  PIN data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 658.280 4.000 658.880 ;
    END
  END data_o[23]
  PIN data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 686.160 4.000 686.760 ;
    END
  END data_o[24]
  PIN data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 714.040 4.000 714.640 ;
    END
  END data_o[25]
  PIN data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 741.920 4.000 742.520 ;
    END
  END data_o[26]
  PIN data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 769.800 4.000 770.400 ;
    END
  END data_o[27]
  PIN data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 797.680 4.000 798.280 ;
    END
  END data_o[28]
  PIN data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 825.560 4.000 826.160 ;
    END
  END data_o[29]
  PIN data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.800 4.000 73.400 ;
    END
  END data_o[2]
  PIN data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 853.440 4.000 854.040 ;
    END
  END data_o[30]
  PIN data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 881.320 4.000 881.920 ;
    END
  END data_o[31]
  PIN data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 4.000 101.280 ;
    END
  END data_o[3]
  PIN data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 128.560 4.000 129.160 ;
    END
  END data_o[4]
  PIN data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END data_o[5]
  PIN data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 184.320 4.000 184.920 ;
    END
  END data_o[6]
  PIN data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.200 4.000 212.800 ;
    END
  END data_o[7]
  PIN data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.080 4.000 240.680 ;
    END
  END data_o[8]
  PIN data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 267.960 4.000 268.560 ;
    END
  END data_o[9]
  PIN done
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 577.850 0.000 578.130 4.000 ;
    END
  END done
  PIN enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.170 0.000 321.450 4.000 ;
    END
  END enable
  PIN mem_opdone
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.510 0.000 449.790 4.000 ;
    END
  END mem_opdone
  PIN mem_operation[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.190 0.000 706.470 4.000 ;
    END
  END mem_operation[0]
  PIN mem_operation[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 834.530 0.000 834.810 4.000 ;
    END
  END mem_operation[1]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.830 0.000 193.110 4.000 ;
    END
  END reset
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 886.960 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 886.960 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 894.240 886.805 ;
      LAYER met1 ;
        RECT 4.670 10.640 895.550 896.540 ;
      LAYER met2 ;
        RECT 4.690 895.720 14.530 896.650 ;
        RECT 15.370 895.720 42.590 896.650 ;
        RECT 43.430 895.720 70.650 896.650 ;
        RECT 71.490 895.720 98.710 896.650 ;
        RECT 99.550 895.720 126.770 896.650 ;
        RECT 127.610 895.720 154.830 896.650 ;
        RECT 155.670 895.720 182.890 896.650 ;
        RECT 183.730 895.720 210.950 896.650 ;
        RECT 211.790 895.720 239.010 896.650 ;
        RECT 239.850 895.720 267.070 896.650 ;
        RECT 267.910 895.720 295.130 896.650 ;
        RECT 295.970 895.720 323.190 896.650 ;
        RECT 324.030 895.720 351.250 896.650 ;
        RECT 352.090 895.720 379.310 896.650 ;
        RECT 380.150 895.720 407.370 896.650 ;
        RECT 408.210 895.720 435.430 896.650 ;
        RECT 436.270 895.720 463.490 896.650 ;
        RECT 464.330 895.720 491.550 896.650 ;
        RECT 492.390 895.720 519.610 896.650 ;
        RECT 520.450 895.720 547.670 896.650 ;
        RECT 548.510 895.720 575.730 896.650 ;
        RECT 576.570 895.720 603.790 896.650 ;
        RECT 604.630 895.720 631.850 896.650 ;
        RECT 632.690 895.720 659.910 896.650 ;
        RECT 660.750 895.720 687.970 896.650 ;
        RECT 688.810 895.720 716.030 896.650 ;
        RECT 716.870 895.720 744.090 896.650 ;
        RECT 744.930 895.720 772.150 896.650 ;
        RECT 772.990 895.720 800.210 896.650 ;
        RECT 801.050 895.720 828.270 896.650 ;
        RECT 829.110 895.720 856.330 896.650 ;
        RECT 857.170 895.720 884.390 896.650 ;
        RECT 885.230 895.720 895.530 896.650 ;
        RECT 4.690 4.280 895.530 895.720 ;
        RECT 4.690 4.000 64.210 4.280 ;
        RECT 65.050 4.000 192.550 4.280 ;
        RECT 193.390 4.000 320.890 4.280 ;
        RECT 321.730 4.000 449.230 4.280 ;
        RECT 450.070 4.000 577.570 4.280 ;
        RECT 578.410 4.000 705.910 4.280 ;
        RECT 706.750 4.000 834.250 4.280 ;
        RECT 835.090 4.000 895.530 4.280 ;
      LAYER met3 ;
        RECT 4.000 882.320 896.000 886.885 ;
        RECT 4.400 880.920 895.600 882.320 ;
        RECT 4.000 854.440 896.000 880.920 ;
        RECT 4.400 853.040 895.600 854.440 ;
        RECT 4.000 826.560 896.000 853.040 ;
        RECT 4.400 825.160 895.600 826.560 ;
        RECT 4.000 798.680 896.000 825.160 ;
        RECT 4.400 797.280 895.600 798.680 ;
        RECT 4.000 770.800 896.000 797.280 ;
        RECT 4.400 769.400 895.600 770.800 ;
        RECT 4.000 742.920 896.000 769.400 ;
        RECT 4.400 741.520 895.600 742.920 ;
        RECT 4.000 715.040 896.000 741.520 ;
        RECT 4.400 713.640 895.600 715.040 ;
        RECT 4.000 687.160 896.000 713.640 ;
        RECT 4.400 685.760 895.600 687.160 ;
        RECT 4.000 659.280 896.000 685.760 ;
        RECT 4.400 657.880 895.600 659.280 ;
        RECT 4.000 631.400 896.000 657.880 ;
        RECT 4.400 630.000 895.600 631.400 ;
        RECT 4.000 603.520 896.000 630.000 ;
        RECT 4.400 602.120 895.600 603.520 ;
        RECT 4.000 575.640 896.000 602.120 ;
        RECT 4.400 574.240 895.600 575.640 ;
        RECT 4.000 547.760 896.000 574.240 ;
        RECT 4.400 546.360 895.600 547.760 ;
        RECT 4.000 519.880 896.000 546.360 ;
        RECT 4.400 518.480 895.600 519.880 ;
        RECT 4.000 492.000 896.000 518.480 ;
        RECT 4.400 490.600 895.600 492.000 ;
        RECT 4.000 464.120 896.000 490.600 ;
        RECT 4.400 462.720 895.600 464.120 ;
        RECT 4.000 436.240 896.000 462.720 ;
        RECT 4.400 434.840 895.600 436.240 ;
        RECT 4.000 408.360 896.000 434.840 ;
        RECT 4.400 406.960 895.600 408.360 ;
        RECT 4.000 380.480 896.000 406.960 ;
        RECT 4.400 379.080 895.600 380.480 ;
        RECT 4.000 352.600 896.000 379.080 ;
        RECT 4.400 351.200 895.600 352.600 ;
        RECT 4.000 324.720 896.000 351.200 ;
        RECT 4.400 323.320 895.600 324.720 ;
        RECT 4.000 296.840 896.000 323.320 ;
        RECT 4.400 295.440 895.600 296.840 ;
        RECT 4.000 268.960 896.000 295.440 ;
        RECT 4.400 267.560 895.600 268.960 ;
        RECT 4.000 241.080 896.000 267.560 ;
        RECT 4.400 239.680 895.600 241.080 ;
        RECT 4.000 213.200 896.000 239.680 ;
        RECT 4.400 211.800 895.600 213.200 ;
        RECT 4.000 185.320 896.000 211.800 ;
        RECT 4.400 183.920 895.600 185.320 ;
        RECT 4.000 157.440 896.000 183.920 ;
        RECT 4.400 156.040 895.600 157.440 ;
        RECT 4.000 129.560 896.000 156.040 ;
        RECT 4.400 128.160 895.600 129.560 ;
        RECT 4.000 101.680 896.000 128.160 ;
        RECT 4.400 100.280 895.600 101.680 ;
        RECT 4.000 73.800 896.000 100.280 ;
        RECT 4.400 72.400 895.600 73.800 ;
        RECT 4.000 45.920 896.000 72.400 ;
        RECT 4.400 44.520 895.600 45.920 ;
        RECT 4.000 18.040 896.000 44.520 ;
        RECT 4.400 16.640 895.600 18.040 ;
        RECT 4.000 10.715 896.000 16.640 ;
      LAYER met4 ;
        RECT 15.015 11.735 20.640 882.465 ;
        RECT 23.040 11.735 97.440 882.465 ;
        RECT 99.840 11.735 174.240 882.465 ;
        RECT 176.640 11.735 251.040 882.465 ;
        RECT 253.440 11.735 327.840 882.465 ;
        RECT 330.240 11.735 404.640 882.465 ;
        RECT 407.040 11.735 481.440 882.465 ;
        RECT 483.840 11.735 558.240 882.465 ;
        RECT 560.640 11.735 635.040 882.465 ;
        RECT 637.440 11.735 711.840 882.465 ;
        RECT 714.240 11.735 788.640 882.465 ;
        RECT 791.040 11.735 825.865 882.465 ;
  END
END Matrix_Multiplication
END LIBRARY

