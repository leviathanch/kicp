version https://git-lfs.github.com/spec/v1
oid sha256:1f8e422422692944a14fad016b92e548c4c0046a94ee8cc8c86a9706f1ce49e8
size 19648
