version https://git-lfs.github.com/spec/v1
oid sha256:31fd30fb74d264b4ce3ee8c4c766689859f3297d239d35e7380fd0c674e407f7
size 165719
