version https://git-lfs.github.com/spec/v1
oid sha256:7984efe386094b56ed877b5cbf9c950be3acbb021ad8b7219201dc1bc3a90973
size 23413
