version https://git-lfs.github.com/spec/v1
oid sha256:1df1b5fb9f965a03353a1afb6942a86073fc96b76a11869f04743d4c80021b22
size 23405
