version https://git-lfs.github.com/spec/v1
oid sha256:c2235a219d097694ba199e6a37d07826a5dce3e26cd039317e520afa1921abb2
size 115943
