magic
tech sky130A
magscale 1 2
timestamp 1685820219
<< nwell >>
rect 1066 176517 178886 177083
rect 1066 175429 178886 175995
rect 1066 174341 178886 174907
rect 1066 173253 178886 173819
rect 1066 172165 178886 172731
rect 1066 171077 178886 171643
rect 1066 169989 178886 170555
rect 1066 168901 178886 169467
rect 1066 167813 178886 168379
rect 1066 166725 178886 167291
rect 1066 165637 178886 166203
rect 1066 164549 178886 165115
rect 1066 163461 178886 164027
rect 1066 162373 178886 162939
rect 1066 161285 178886 161851
rect 1066 160197 178886 160763
rect 1066 159109 178886 159675
rect 1066 158021 178886 158587
rect 1066 156933 178886 157499
rect 1066 155845 178886 156411
rect 1066 154757 178886 155323
rect 1066 153669 178886 154235
rect 1066 152581 178886 153147
rect 1066 151493 178886 152059
rect 1066 150405 178886 150971
rect 1066 149317 178886 149883
rect 1066 148229 178886 148795
rect 1066 147141 178886 147707
rect 1066 146053 178886 146619
rect 1066 144965 178886 145531
rect 1066 143877 178886 144443
rect 1066 142789 178886 143355
rect 1066 141701 178886 142267
rect 1066 140613 178886 141179
rect 1066 139525 178886 140091
rect 1066 138437 178886 139003
rect 1066 137349 178886 137915
rect 1066 136261 178886 136827
rect 1066 135173 178886 135739
rect 1066 134085 178886 134651
rect 1066 132997 178886 133563
rect 1066 131909 178886 132475
rect 1066 130821 178886 131387
rect 1066 129733 178886 130299
rect 1066 128645 178886 129211
rect 1066 127557 178886 128123
rect 1066 126469 178886 127035
rect 1066 125381 178886 125947
rect 1066 124293 178886 124859
rect 1066 123205 178886 123771
rect 1066 122117 178886 122683
rect 1066 121029 178886 121595
rect 1066 119941 178886 120507
rect 1066 118853 178886 119419
rect 1066 117765 178886 118331
rect 1066 116677 178886 117243
rect 1066 115589 178886 116155
rect 1066 114501 178886 115067
rect 1066 113413 178886 113979
rect 1066 112325 178886 112891
rect 1066 111237 178886 111803
rect 1066 110149 178886 110715
rect 1066 109061 178886 109627
rect 1066 107973 178886 108539
rect 1066 106885 178886 107451
rect 1066 105797 178886 106363
rect 1066 104709 178886 105275
rect 1066 103621 178886 104187
rect 1066 102533 178886 103099
rect 1066 101445 178886 102011
rect 1066 100357 178886 100923
rect 1066 99269 178886 99835
rect 1066 98181 178886 98747
rect 1066 97093 178886 97659
rect 1066 96005 178886 96571
rect 1066 94917 178886 95483
rect 1066 93829 178886 94395
rect 1066 92741 178886 93307
rect 1066 91653 178886 92219
rect 1066 90565 178886 91131
rect 1066 89477 178886 90043
rect 1066 88389 178886 88955
rect 1066 87301 178886 87867
rect 1066 86213 178886 86779
rect 1066 85125 178886 85691
rect 1066 84037 178886 84603
rect 1066 82949 178886 83515
rect 1066 81861 178886 82427
rect 1066 80773 178886 81339
rect 1066 79685 178886 80251
rect 1066 78597 178886 79163
rect 1066 77509 178886 78075
rect 1066 76421 178886 76987
rect 1066 75333 178886 75899
rect 1066 74245 178886 74811
rect 1066 73157 178886 73723
rect 1066 72069 178886 72635
rect 1066 70981 178886 71547
rect 1066 69893 178886 70459
rect 1066 68805 178886 69371
rect 1066 67717 178886 68283
rect 1066 66629 178886 67195
rect 1066 65541 178886 66107
rect 1066 64453 178886 65019
rect 1066 63365 178886 63931
rect 1066 62277 178886 62843
rect 1066 61189 178886 61755
rect 1066 60101 178886 60667
rect 1066 59013 178886 59579
rect 1066 57925 178886 58491
rect 1066 56837 178886 57403
rect 1066 55749 178886 56315
rect 1066 54661 178886 55227
rect 1066 53573 178886 54139
rect 1066 52485 178886 53051
rect 1066 51397 178886 51963
rect 1066 50309 178886 50875
rect 1066 49221 178886 49787
rect 1066 48133 178886 48699
rect 1066 47045 178886 47611
rect 1066 45957 178886 46523
rect 1066 44869 178886 45435
rect 1066 43781 178886 44347
rect 1066 42693 178886 43259
rect 1066 41605 178886 42171
rect 1066 40517 178886 41083
rect 1066 39429 178886 39995
rect 1066 38341 178886 38907
rect 1066 37253 178886 37819
rect 1066 36165 178886 36731
rect 1066 35077 178886 35643
rect 1066 33989 178886 34555
rect 1066 32901 178886 33467
rect 1066 31813 178886 32379
rect 1066 30725 178886 31291
rect 1066 29637 178886 30203
rect 1066 28549 178886 29115
rect 1066 27461 178886 28027
rect 1066 26373 178886 26939
rect 1066 25285 178886 25851
rect 1066 24197 178886 24763
rect 1066 23109 178886 23675
rect 1066 22021 178886 22587
rect 1066 20933 178886 21499
rect 1066 19845 178886 20411
rect 1066 18757 178886 19323
rect 1066 17669 178886 18235
rect 1066 16581 178886 17147
rect 1066 15493 178886 16059
rect 1066 14405 178886 14971
rect 1066 13317 178886 13883
rect 1066 12229 178886 12795
rect 1066 11141 178886 11707
rect 1066 10053 178886 10619
rect 1066 8965 178886 9531
rect 1066 7877 178886 8443
rect 1066 6789 178886 7355
rect 1066 5701 178886 6267
rect 1066 4613 178886 5179
rect 1066 3525 178886 4091
rect 1066 2437 178886 3003
<< obsli1 >>
rect 1104 2159 178848 177361
<< obsm1 >>
rect 1104 76 178848 177392
<< metal2 >>
rect 5446 0 5502 800
rect 7102 0 7158 800
rect 8758 0 8814 800
rect 10414 0 10470 800
rect 12070 0 12126 800
rect 13726 0 13782 800
rect 15382 0 15438 800
rect 17038 0 17094 800
rect 18694 0 18750 800
rect 20350 0 20406 800
rect 22006 0 22062 800
rect 23662 0 23718 800
rect 25318 0 25374 800
rect 26974 0 27030 800
rect 28630 0 28686 800
rect 30286 0 30342 800
rect 31942 0 31998 800
rect 33598 0 33654 800
rect 35254 0 35310 800
rect 36910 0 36966 800
rect 38566 0 38622 800
rect 40222 0 40278 800
rect 41878 0 41934 800
rect 43534 0 43590 800
rect 45190 0 45246 800
rect 46846 0 46902 800
rect 48502 0 48558 800
rect 50158 0 50214 800
rect 51814 0 51870 800
rect 53470 0 53526 800
rect 55126 0 55182 800
rect 56782 0 56838 800
rect 58438 0 58494 800
rect 60094 0 60150 800
rect 61750 0 61806 800
rect 63406 0 63462 800
rect 65062 0 65118 800
rect 66718 0 66774 800
rect 68374 0 68430 800
rect 70030 0 70086 800
rect 71686 0 71742 800
rect 73342 0 73398 800
rect 74998 0 75054 800
rect 76654 0 76710 800
rect 78310 0 78366 800
rect 79966 0 80022 800
rect 81622 0 81678 800
rect 83278 0 83334 800
rect 84934 0 84990 800
rect 86590 0 86646 800
rect 88246 0 88302 800
rect 89902 0 89958 800
rect 91558 0 91614 800
rect 93214 0 93270 800
rect 94870 0 94926 800
rect 96526 0 96582 800
rect 98182 0 98238 800
rect 99838 0 99894 800
rect 101494 0 101550 800
rect 103150 0 103206 800
rect 104806 0 104862 800
rect 106462 0 106518 800
rect 108118 0 108174 800
rect 109774 0 109830 800
rect 111430 0 111486 800
rect 113086 0 113142 800
rect 114742 0 114798 800
rect 116398 0 116454 800
rect 118054 0 118110 800
rect 119710 0 119766 800
rect 121366 0 121422 800
rect 123022 0 123078 800
rect 124678 0 124734 800
rect 126334 0 126390 800
rect 127990 0 128046 800
rect 129646 0 129702 800
rect 131302 0 131358 800
rect 132958 0 133014 800
rect 134614 0 134670 800
rect 136270 0 136326 800
rect 137926 0 137982 800
rect 139582 0 139638 800
rect 141238 0 141294 800
rect 142894 0 142950 800
rect 144550 0 144606 800
rect 146206 0 146262 800
rect 147862 0 147918 800
rect 149518 0 149574 800
rect 151174 0 151230 800
rect 152830 0 152886 800
rect 154486 0 154542 800
rect 156142 0 156198 800
rect 157798 0 157854 800
rect 159454 0 159510 800
rect 161110 0 161166 800
rect 162766 0 162822 800
rect 164422 0 164478 800
rect 166078 0 166134 800
rect 167734 0 167790 800
rect 169390 0 169446 800
rect 171046 0 171102 800
rect 172702 0 172758 800
rect 174358 0 174414 800
<< obsm2 >>
rect 1584 856 178368 177381
rect 1584 31 5390 856
rect 5558 31 7046 856
rect 7214 31 8702 856
rect 8870 31 10358 856
rect 10526 31 12014 856
rect 12182 31 13670 856
rect 13838 31 15326 856
rect 15494 31 16982 856
rect 17150 31 18638 856
rect 18806 31 20294 856
rect 20462 31 21950 856
rect 22118 31 23606 856
rect 23774 31 25262 856
rect 25430 31 26918 856
rect 27086 31 28574 856
rect 28742 31 30230 856
rect 30398 31 31886 856
rect 32054 31 33542 856
rect 33710 31 35198 856
rect 35366 31 36854 856
rect 37022 31 38510 856
rect 38678 31 40166 856
rect 40334 31 41822 856
rect 41990 31 43478 856
rect 43646 31 45134 856
rect 45302 31 46790 856
rect 46958 31 48446 856
rect 48614 31 50102 856
rect 50270 31 51758 856
rect 51926 31 53414 856
rect 53582 31 55070 856
rect 55238 31 56726 856
rect 56894 31 58382 856
rect 58550 31 60038 856
rect 60206 31 61694 856
rect 61862 31 63350 856
rect 63518 31 65006 856
rect 65174 31 66662 856
rect 66830 31 68318 856
rect 68486 31 69974 856
rect 70142 31 71630 856
rect 71798 31 73286 856
rect 73454 31 74942 856
rect 75110 31 76598 856
rect 76766 31 78254 856
rect 78422 31 79910 856
rect 80078 31 81566 856
rect 81734 31 83222 856
rect 83390 31 84878 856
rect 85046 31 86534 856
rect 86702 31 88190 856
rect 88358 31 89846 856
rect 90014 31 91502 856
rect 91670 31 93158 856
rect 93326 31 94814 856
rect 94982 31 96470 856
rect 96638 31 98126 856
rect 98294 31 99782 856
rect 99950 31 101438 856
rect 101606 31 103094 856
rect 103262 31 104750 856
rect 104918 31 106406 856
rect 106574 31 108062 856
rect 108230 31 109718 856
rect 109886 31 111374 856
rect 111542 31 113030 856
rect 113198 31 114686 856
rect 114854 31 116342 856
rect 116510 31 117998 856
rect 118166 31 119654 856
rect 119822 31 121310 856
rect 121478 31 122966 856
rect 123134 31 124622 856
rect 124790 31 126278 856
rect 126446 31 127934 856
rect 128102 31 129590 856
rect 129758 31 131246 856
rect 131414 31 132902 856
rect 133070 31 134558 856
rect 134726 31 136214 856
rect 136382 31 137870 856
rect 138038 31 139526 856
rect 139694 31 141182 856
rect 141350 31 142838 856
rect 143006 31 144494 856
rect 144662 31 146150 856
rect 146318 31 147806 856
rect 147974 31 149462 856
rect 149630 31 151118 856
rect 151286 31 152774 856
rect 152942 31 154430 856
rect 154598 31 156086 856
rect 156254 31 157742 856
rect 157910 31 159398 856
rect 159566 31 161054 856
rect 161222 31 162710 856
rect 162878 31 164366 856
rect 164534 31 166022 856
rect 166190 31 167678 856
rect 167846 31 169334 856
rect 169502 31 170990 856
rect 171158 31 172646 856
rect 172814 31 174302 856
rect 174470 31 178368 856
<< obsm3 >>
rect 2681 35 178283 177377
<< metal4 >>
rect 4208 2128 4528 177392
rect 19568 2128 19888 177392
rect 34928 2128 35248 177392
rect 50288 2128 50608 177392
rect 65648 2128 65968 177392
rect 81008 2128 81328 177392
rect 96368 2128 96688 177392
rect 111728 2128 112048 177392
rect 127088 2128 127408 177392
rect 142448 2128 142768 177392
rect 157808 2128 158128 177392
rect 173168 2128 173488 177392
<< obsm4 >>
rect 3003 2048 4128 154053
rect 4608 2048 19488 154053
rect 19968 2048 34848 154053
rect 35328 2048 50208 154053
rect 50688 2048 65568 154053
rect 66048 2048 80928 154053
rect 81408 2048 96288 154053
rect 96768 2048 111648 154053
rect 112128 2048 127008 154053
rect 127488 2048 142368 154053
rect 142848 2048 157728 154053
rect 158208 2048 173088 154053
rect 173568 2048 175661 154053
rect 3003 35 175661 2048
<< labels >>
rlabel metal2 s 13726 0 13782 800 6 addr_o[0]
port 1 nsew signal output
rlabel metal2 s 66718 0 66774 800 6 addr_o[10]
port 2 nsew signal output
rlabel metal2 s 71686 0 71742 800 6 addr_o[11]
port 3 nsew signal output
rlabel metal2 s 76654 0 76710 800 6 addr_o[12]
port 4 nsew signal output
rlabel metal2 s 81622 0 81678 800 6 addr_o[13]
port 5 nsew signal output
rlabel metal2 s 86590 0 86646 800 6 addr_o[14]
port 6 nsew signal output
rlabel metal2 s 91558 0 91614 800 6 addr_o[15]
port 7 nsew signal output
rlabel metal2 s 96526 0 96582 800 6 addr_o[16]
port 8 nsew signal output
rlabel metal2 s 101494 0 101550 800 6 addr_o[17]
port 9 nsew signal output
rlabel metal2 s 106462 0 106518 800 6 addr_o[18]
port 10 nsew signal output
rlabel metal2 s 111430 0 111486 800 6 addr_o[19]
port 11 nsew signal output
rlabel metal2 s 20350 0 20406 800 6 addr_o[1]
port 12 nsew signal output
rlabel metal2 s 116398 0 116454 800 6 addr_o[20]
port 13 nsew signal output
rlabel metal2 s 121366 0 121422 800 6 addr_o[21]
port 14 nsew signal output
rlabel metal2 s 126334 0 126390 800 6 addr_o[22]
port 15 nsew signal output
rlabel metal2 s 131302 0 131358 800 6 addr_o[23]
port 16 nsew signal output
rlabel metal2 s 136270 0 136326 800 6 addr_o[24]
port 17 nsew signal output
rlabel metal2 s 141238 0 141294 800 6 addr_o[25]
port 18 nsew signal output
rlabel metal2 s 146206 0 146262 800 6 addr_o[26]
port 19 nsew signal output
rlabel metal2 s 151174 0 151230 800 6 addr_o[27]
port 20 nsew signal output
rlabel metal2 s 156142 0 156198 800 6 addr_o[28]
port 21 nsew signal output
rlabel metal2 s 161110 0 161166 800 6 addr_o[29]
port 22 nsew signal output
rlabel metal2 s 26974 0 27030 800 6 addr_o[2]
port 23 nsew signal output
rlabel metal2 s 166078 0 166134 800 6 addr_o[30]
port 24 nsew signal output
rlabel metal2 s 171046 0 171102 800 6 addr_o[31]
port 25 nsew signal output
rlabel metal2 s 31942 0 31998 800 6 addr_o[3]
port 26 nsew signal output
rlabel metal2 s 36910 0 36966 800 6 addr_o[4]
port 27 nsew signal output
rlabel metal2 s 41878 0 41934 800 6 addr_o[5]
port 28 nsew signal output
rlabel metal2 s 46846 0 46902 800 6 addr_o[6]
port 29 nsew signal output
rlabel metal2 s 51814 0 51870 800 6 addr_o[7]
port 30 nsew signal output
rlabel metal2 s 56782 0 56838 800 6 addr_o[8]
port 31 nsew signal output
rlabel metal2 s 61750 0 61806 800 6 addr_o[9]
port 32 nsew signal output
rlabel metal2 s 5446 0 5502 800 6 clk
port 33 nsew signal input
rlabel metal2 s 15382 0 15438 800 6 data_i[0]
port 34 nsew signal input
rlabel metal2 s 68374 0 68430 800 6 data_i[10]
port 35 nsew signal input
rlabel metal2 s 73342 0 73398 800 6 data_i[11]
port 36 nsew signal input
rlabel metal2 s 78310 0 78366 800 6 data_i[12]
port 37 nsew signal input
rlabel metal2 s 83278 0 83334 800 6 data_i[13]
port 38 nsew signal input
rlabel metal2 s 88246 0 88302 800 6 data_i[14]
port 39 nsew signal input
rlabel metal2 s 93214 0 93270 800 6 data_i[15]
port 40 nsew signal input
rlabel metal2 s 98182 0 98238 800 6 data_i[16]
port 41 nsew signal input
rlabel metal2 s 103150 0 103206 800 6 data_i[17]
port 42 nsew signal input
rlabel metal2 s 108118 0 108174 800 6 data_i[18]
port 43 nsew signal input
rlabel metal2 s 113086 0 113142 800 6 data_i[19]
port 44 nsew signal input
rlabel metal2 s 22006 0 22062 800 6 data_i[1]
port 45 nsew signal input
rlabel metal2 s 118054 0 118110 800 6 data_i[20]
port 46 nsew signal input
rlabel metal2 s 123022 0 123078 800 6 data_i[21]
port 47 nsew signal input
rlabel metal2 s 127990 0 128046 800 6 data_i[22]
port 48 nsew signal input
rlabel metal2 s 132958 0 133014 800 6 data_i[23]
port 49 nsew signal input
rlabel metal2 s 137926 0 137982 800 6 data_i[24]
port 50 nsew signal input
rlabel metal2 s 142894 0 142950 800 6 data_i[25]
port 51 nsew signal input
rlabel metal2 s 147862 0 147918 800 6 data_i[26]
port 52 nsew signal input
rlabel metal2 s 152830 0 152886 800 6 data_i[27]
port 53 nsew signal input
rlabel metal2 s 157798 0 157854 800 6 data_i[28]
port 54 nsew signal input
rlabel metal2 s 162766 0 162822 800 6 data_i[29]
port 55 nsew signal input
rlabel metal2 s 28630 0 28686 800 6 data_i[2]
port 56 nsew signal input
rlabel metal2 s 167734 0 167790 800 6 data_i[30]
port 57 nsew signal input
rlabel metal2 s 172702 0 172758 800 6 data_i[31]
port 58 nsew signal input
rlabel metal2 s 33598 0 33654 800 6 data_i[3]
port 59 nsew signal input
rlabel metal2 s 38566 0 38622 800 6 data_i[4]
port 60 nsew signal input
rlabel metal2 s 43534 0 43590 800 6 data_i[5]
port 61 nsew signal input
rlabel metal2 s 48502 0 48558 800 6 data_i[6]
port 62 nsew signal input
rlabel metal2 s 53470 0 53526 800 6 data_i[7]
port 63 nsew signal input
rlabel metal2 s 58438 0 58494 800 6 data_i[8]
port 64 nsew signal input
rlabel metal2 s 63406 0 63462 800 6 data_i[9]
port 65 nsew signal input
rlabel metal2 s 17038 0 17094 800 6 data_o[0]
port 66 nsew signal output
rlabel metal2 s 70030 0 70086 800 6 data_o[10]
port 67 nsew signal output
rlabel metal2 s 74998 0 75054 800 6 data_o[11]
port 68 nsew signal output
rlabel metal2 s 79966 0 80022 800 6 data_o[12]
port 69 nsew signal output
rlabel metal2 s 84934 0 84990 800 6 data_o[13]
port 70 nsew signal output
rlabel metal2 s 89902 0 89958 800 6 data_o[14]
port 71 nsew signal output
rlabel metal2 s 94870 0 94926 800 6 data_o[15]
port 72 nsew signal output
rlabel metal2 s 99838 0 99894 800 6 data_o[16]
port 73 nsew signal output
rlabel metal2 s 104806 0 104862 800 6 data_o[17]
port 74 nsew signal output
rlabel metal2 s 109774 0 109830 800 6 data_o[18]
port 75 nsew signal output
rlabel metal2 s 114742 0 114798 800 6 data_o[19]
port 76 nsew signal output
rlabel metal2 s 23662 0 23718 800 6 data_o[1]
port 77 nsew signal output
rlabel metal2 s 119710 0 119766 800 6 data_o[20]
port 78 nsew signal output
rlabel metal2 s 124678 0 124734 800 6 data_o[21]
port 79 nsew signal output
rlabel metal2 s 129646 0 129702 800 6 data_o[22]
port 80 nsew signal output
rlabel metal2 s 134614 0 134670 800 6 data_o[23]
port 81 nsew signal output
rlabel metal2 s 139582 0 139638 800 6 data_o[24]
port 82 nsew signal output
rlabel metal2 s 144550 0 144606 800 6 data_o[25]
port 83 nsew signal output
rlabel metal2 s 149518 0 149574 800 6 data_o[26]
port 84 nsew signal output
rlabel metal2 s 154486 0 154542 800 6 data_o[27]
port 85 nsew signal output
rlabel metal2 s 159454 0 159510 800 6 data_o[28]
port 86 nsew signal output
rlabel metal2 s 164422 0 164478 800 6 data_o[29]
port 87 nsew signal output
rlabel metal2 s 30286 0 30342 800 6 data_o[2]
port 88 nsew signal output
rlabel metal2 s 169390 0 169446 800 6 data_o[30]
port 89 nsew signal output
rlabel metal2 s 174358 0 174414 800 6 data_o[31]
port 90 nsew signal output
rlabel metal2 s 35254 0 35310 800 6 data_o[3]
port 91 nsew signal output
rlabel metal2 s 40222 0 40278 800 6 data_o[4]
port 92 nsew signal output
rlabel metal2 s 45190 0 45246 800 6 data_o[5]
port 93 nsew signal output
rlabel metal2 s 50158 0 50214 800 6 data_o[6]
port 94 nsew signal output
rlabel metal2 s 55126 0 55182 800 6 data_o[7]
port 95 nsew signal output
rlabel metal2 s 60094 0 60150 800 6 data_o[8]
port 96 nsew signal output
rlabel metal2 s 65062 0 65118 800 6 data_o[9]
port 97 nsew signal output
rlabel metal2 s 12070 0 12126 800 6 done
port 98 nsew signal output
rlabel metal2 s 8758 0 8814 800 6 enable
port 99 nsew signal input
rlabel metal2 s 10414 0 10470 800 6 mem_opdone
port 100 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 mem_operation[0]
port 101 nsew signal output
rlabel metal2 s 25318 0 25374 800 6 mem_operation[1]
port 102 nsew signal output
rlabel metal2 s 7102 0 7158 800 6 reset
port 103 nsew signal input
rlabel metal4 s 4208 2128 4528 177392 6 vccd1
port 104 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 177392 6 vccd1
port 104 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 177392 6 vccd1
port 104 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 177392 6 vccd1
port 104 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 177392 6 vccd1
port 104 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 177392 6 vccd1
port 104 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 177392 6 vssd1
port 105 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 177392 6 vssd1
port 105 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 177392 6 vssd1
port 105 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 177392 6 vssd1
port 105 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 177392 6 vssd1
port 105 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 177392 6 vssd1
port 105 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 180000 180000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 61415790
string GDS_FILE /home/leviathan/kicp/openlane/Matrix_Convolution/runs/23_06_03_19_10/results/signoff/Matrix_Convolution.magic.gds
string GDS_START 1560760
<< end >>

