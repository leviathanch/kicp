magic
tech sky130A
magscale 1 2
timestamp 1685822584
<< obsli1 >>
rect 1104 2159 498824 297585
<< obsm1 >>
rect 934 76 499086 297616
<< metal2 >>
rect 2502 0 2558 800
rect 3514 0 3570 800
rect 4526 0 4582 800
rect 5538 0 5594 800
rect 6550 0 6606 800
rect 7562 0 7618 800
rect 8574 0 8630 800
rect 9586 0 9642 800
rect 10598 0 10654 800
rect 11610 0 11666 800
rect 12622 0 12678 800
rect 13634 0 13690 800
rect 14646 0 14702 800
rect 15658 0 15714 800
rect 16670 0 16726 800
rect 17682 0 17738 800
rect 18694 0 18750 800
rect 19706 0 19762 800
rect 20718 0 20774 800
rect 21730 0 21786 800
rect 22742 0 22798 800
rect 23754 0 23810 800
rect 24766 0 24822 800
rect 25778 0 25834 800
rect 26790 0 26846 800
rect 27802 0 27858 800
rect 28814 0 28870 800
rect 29826 0 29882 800
rect 30838 0 30894 800
rect 31850 0 31906 800
rect 32862 0 32918 800
rect 33874 0 33930 800
rect 34886 0 34942 800
rect 35898 0 35954 800
rect 36910 0 36966 800
rect 37922 0 37978 800
rect 38934 0 38990 800
rect 39946 0 40002 800
rect 40958 0 41014 800
rect 41970 0 42026 800
rect 42982 0 43038 800
rect 43994 0 44050 800
rect 45006 0 45062 800
rect 46018 0 46074 800
rect 47030 0 47086 800
rect 48042 0 48098 800
rect 49054 0 49110 800
rect 50066 0 50122 800
rect 51078 0 51134 800
rect 52090 0 52146 800
rect 53102 0 53158 800
rect 54114 0 54170 800
rect 55126 0 55182 800
rect 56138 0 56194 800
rect 57150 0 57206 800
rect 58162 0 58218 800
rect 59174 0 59230 800
rect 60186 0 60242 800
rect 61198 0 61254 800
rect 62210 0 62266 800
rect 63222 0 63278 800
rect 64234 0 64290 800
rect 65246 0 65302 800
rect 66258 0 66314 800
rect 67270 0 67326 800
rect 68282 0 68338 800
rect 69294 0 69350 800
rect 70306 0 70362 800
rect 71318 0 71374 800
rect 72330 0 72386 800
rect 73342 0 73398 800
rect 74354 0 74410 800
rect 75366 0 75422 800
rect 76378 0 76434 800
rect 77390 0 77446 800
rect 78402 0 78458 800
rect 79414 0 79470 800
rect 80426 0 80482 800
rect 81438 0 81494 800
rect 82450 0 82506 800
rect 83462 0 83518 800
rect 84474 0 84530 800
rect 85486 0 85542 800
rect 86498 0 86554 800
rect 87510 0 87566 800
rect 88522 0 88578 800
rect 89534 0 89590 800
rect 90546 0 90602 800
rect 91558 0 91614 800
rect 92570 0 92626 800
rect 93582 0 93638 800
rect 94594 0 94650 800
rect 95606 0 95662 800
rect 96618 0 96674 800
rect 97630 0 97686 800
rect 98642 0 98698 800
rect 99654 0 99710 800
rect 100666 0 100722 800
rect 101678 0 101734 800
rect 102690 0 102746 800
rect 103702 0 103758 800
rect 104714 0 104770 800
rect 105726 0 105782 800
rect 106738 0 106794 800
rect 107750 0 107806 800
rect 108762 0 108818 800
rect 109774 0 109830 800
rect 110786 0 110842 800
rect 111798 0 111854 800
rect 112810 0 112866 800
rect 113822 0 113878 800
rect 114834 0 114890 800
rect 115846 0 115902 800
rect 116858 0 116914 800
rect 117870 0 117926 800
rect 118882 0 118938 800
rect 119894 0 119950 800
rect 120906 0 120962 800
rect 121918 0 121974 800
rect 122930 0 122986 800
rect 123942 0 123998 800
rect 124954 0 125010 800
rect 125966 0 126022 800
rect 126978 0 127034 800
rect 127990 0 128046 800
rect 129002 0 129058 800
rect 130014 0 130070 800
rect 131026 0 131082 800
rect 132038 0 132094 800
rect 133050 0 133106 800
rect 134062 0 134118 800
rect 135074 0 135130 800
rect 136086 0 136142 800
rect 137098 0 137154 800
rect 138110 0 138166 800
rect 139122 0 139178 800
rect 140134 0 140190 800
rect 141146 0 141202 800
rect 142158 0 142214 800
rect 143170 0 143226 800
rect 144182 0 144238 800
rect 145194 0 145250 800
rect 146206 0 146262 800
rect 147218 0 147274 800
rect 148230 0 148286 800
rect 149242 0 149298 800
rect 150254 0 150310 800
rect 151266 0 151322 800
rect 152278 0 152334 800
rect 153290 0 153346 800
rect 154302 0 154358 800
rect 155314 0 155370 800
rect 156326 0 156382 800
rect 157338 0 157394 800
rect 158350 0 158406 800
rect 159362 0 159418 800
rect 160374 0 160430 800
rect 161386 0 161442 800
rect 162398 0 162454 800
rect 163410 0 163466 800
rect 164422 0 164478 800
rect 165434 0 165490 800
rect 166446 0 166502 800
rect 167458 0 167514 800
rect 168470 0 168526 800
rect 169482 0 169538 800
rect 170494 0 170550 800
rect 171506 0 171562 800
rect 172518 0 172574 800
rect 173530 0 173586 800
rect 174542 0 174598 800
rect 175554 0 175610 800
rect 176566 0 176622 800
rect 177578 0 177634 800
rect 178590 0 178646 800
rect 179602 0 179658 800
rect 180614 0 180670 800
rect 181626 0 181682 800
rect 182638 0 182694 800
rect 183650 0 183706 800
rect 184662 0 184718 800
rect 185674 0 185730 800
rect 186686 0 186742 800
rect 187698 0 187754 800
rect 188710 0 188766 800
rect 189722 0 189778 800
rect 190734 0 190790 800
rect 191746 0 191802 800
rect 192758 0 192814 800
rect 193770 0 193826 800
rect 194782 0 194838 800
rect 195794 0 195850 800
rect 196806 0 196862 800
rect 197818 0 197874 800
rect 198830 0 198886 800
rect 199842 0 199898 800
rect 200854 0 200910 800
rect 201866 0 201922 800
rect 202878 0 202934 800
rect 203890 0 203946 800
rect 204902 0 204958 800
rect 205914 0 205970 800
rect 206926 0 206982 800
rect 207938 0 207994 800
rect 208950 0 209006 800
rect 209962 0 210018 800
rect 210974 0 211030 800
rect 211986 0 212042 800
rect 212998 0 213054 800
rect 214010 0 214066 800
rect 215022 0 215078 800
rect 216034 0 216090 800
rect 217046 0 217102 800
rect 218058 0 218114 800
rect 219070 0 219126 800
rect 220082 0 220138 800
rect 221094 0 221150 800
rect 222106 0 222162 800
rect 223118 0 223174 800
rect 224130 0 224186 800
rect 225142 0 225198 800
rect 226154 0 226210 800
rect 227166 0 227222 800
rect 228178 0 228234 800
rect 229190 0 229246 800
rect 230202 0 230258 800
rect 231214 0 231270 800
rect 232226 0 232282 800
rect 233238 0 233294 800
rect 234250 0 234306 800
rect 235262 0 235318 800
rect 236274 0 236330 800
rect 237286 0 237342 800
rect 238298 0 238354 800
rect 239310 0 239366 800
rect 240322 0 240378 800
rect 241334 0 241390 800
rect 242346 0 242402 800
rect 243358 0 243414 800
rect 244370 0 244426 800
rect 245382 0 245438 800
rect 246394 0 246450 800
rect 247406 0 247462 800
rect 248418 0 248474 800
rect 249430 0 249486 800
rect 250442 0 250498 800
rect 251454 0 251510 800
rect 252466 0 252522 800
rect 253478 0 253534 800
rect 254490 0 254546 800
rect 255502 0 255558 800
rect 256514 0 256570 800
rect 257526 0 257582 800
rect 258538 0 258594 800
rect 259550 0 259606 800
rect 260562 0 260618 800
rect 261574 0 261630 800
rect 262586 0 262642 800
rect 263598 0 263654 800
rect 264610 0 264666 800
rect 265622 0 265678 800
rect 266634 0 266690 800
rect 267646 0 267702 800
rect 268658 0 268714 800
rect 269670 0 269726 800
rect 270682 0 270738 800
rect 271694 0 271750 800
rect 272706 0 272762 800
rect 273718 0 273774 800
rect 274730 0 274786 800
rect 275742 0 275798 800
rect 276754 0 276810 800
rect 277766 0 277822 800
rect 278778 0 278834 800
rect 279790 0 279846 800
rect 280802 0 280858 800
rect 281814 0 281870 800
rect 282826 0 282882 800
rect 283838 0 283894 800
rect 284850 0 284906 800
rect 285862 0 285918 800
rect 286874 0 286930 800
rect 287886 0 287942 800
rect 288898 0 288954 800
rect 289910 0 289966 800
rect 290922 0 290978 800
rect 291934 0 291990 800
rect 292946 0 293002 800
rect 293958 0 294014 800
rect 294970 0 295026 800
rect 295982 0 296038 800
rect 296994 0 297050 800
rect 298006 0 298062 800
rect 299018 0 299074 800
rect 300030 0 300086 800
rect 301042 0 301098 800
rect 302054 0 302110 800
rect 303066 0 303122 800
rect 304078 0 304134 800
rect 305090 0 305146 800
rect 306102 0 306158 800
rect 307114 0 307170 800
rect 308126 0 308182 800
rect 309138 0 309194 800
rect 310150 0 310206 800
rect 311162 0 311218 800
rect 312174 0 312230 800
rect 313186 0 313242 800
rect 314198 0 314254 800
rect 315210 0 315266 800
rect 316222 0 316278 800
rect 317234 0 317290 800
rect 318246 0 318302 800
rect 319258 0 319314 800
rect 320270 0 320326 800
rect 321282 0 321338 800
rect 322294 0 322350 800
rect 323306 0 323362 800
rect 324318 0 324374 800
rect 325330 0 325386 800
rect 326342 0 326398 800
rect 327354 0 327410 800
rect 328366 0 328422 800
rect 329378 0 329434 800
rect 330390 0 330446 800
rect 331402 0 331458 800
rect 332414 0 332470 800
rect 333426 0 333482 800
rect 334438 0 334494 800
rect 335450 0 335506 800
rect 336462 0 336518 800
rect 337474 0 337530 800
rect 338486 0 338542 800
rect 339498 0 339554 800
rect 340510 0 340566 800
rect 341522 0 341578 800
rect 342534 0 342590 800
rect 343546 0 343602 800
rect 344558 0 344614 800
rect 345570 0 345626 800
rect 346582 0 346638 800
rect 347594 0 347650 800
rect 348606 0 348662 800
rect 349618 0 349674 800
rect 350630 0 350686 800
rect 351642 0 351698 800
rect 352654 0 352710 800
rect 353666 0 353722 800
rect 354678 0 354734 800
rect 355690 0 355746 800
rect 356702 0 356758 800
rect 357714 0 357770 800
rect 358726 0 358782 800
rect 359738 0 359794 800
rect 360750 0 360806 800
rect 361762 0 361818 800
rect 362774 0 362830 800
rect 363786 0 363842 800
rect 364798 0 364854 800
rect 365810 0 365866 800
rect 366822 0 366878 800
rect 367834 0 367890 800
rect 368846 0 368902 800
rect 369858 0 369914 800
rect 370870 0 370926 800
rect 371882 0 371938 800
rect 372894 0 372950 800
rect 373906 0 373962 800
rect 374918 0 374974 800
rect 375930 0 375986 800
rect 376942 0 376998 800
rect 377954 0 378010 800
rect 378966 0 379022 800
rect 379978 0 380034 800
rect 380990 0 381046 800
rect 382002 0 382058 800
rect 383014 0 383070 800
rect 384026 0 384082 800
rect 385038 0 385094 800
rect 386050 0 386106 800
rect 387062 0 387118 800
rect 388074 0 388130 800
rect 389086 0 389142 800
rect 390098 0 390154 800
rect 391110 0 391166 800
rect 392122 0 392178 800
rect 393134 0 393190 800
rect 394146 0 394202 800
rect 395158 0 395214 800
rect 396170 0 396226 800
rect 397182 0 397238 800
rect 398194 0 398250 800
rect 399206 0 399262 800
rect 400218 0 400274 800
rect 401230 0 401286 800
rect 402242 0 402298 800
rect 403254 0 403310 800
rect 404266 0 404322 800
rect 405278 0 405334 800
rect 406290 0 406346 800
rect 407302 0 407358 800
rect 408314 0 408370 800
rect 409326 0 409382 800
rect 410338 0 410394 800
rect 411350 0 411406 800
rect 412362 0 412418 800
rect 413374 0 413430 800
rect 414386 0 414442 800
rect 415398 0 415454 800
rect 416410 0 416466 800
rect 417422 0 417478 800
rect 418434 0 418490 800
rect 419446 0 419502 800
rect 420458 0 420514 800
rect 421470 0 421526 800
rect 422482 0 422538 800
rect 423494 0 423550 800
rect 424506 0 424562 800
rect 425518 0 425574 800
rect 426530 0 426586 800
rect 427542 0 427598 800
rect 428554 0 428610 800
rect 429566 0 429622 800
rect 430578 0 430634 800
rect 431590 0 431646 800
rect 432602 0 432658 800
rect 433614 0 433670 800
rect 434626 0 434682 800
rect 435638 0 435694 800
rect 436650 0 436706 800
rect 437662 0 437718 800
rect 438674 0 438730 800
rect 439686 0 439742 800
rect 440698 0 440754 800
rect 441710 0 441766 800
rect 442722 0 442778 800
rect 443734 0 443790 800
rect 444746 0 444802 800
rect 445758 0 445814 800
rect 446770 0 446826 800
rect 447782 0 447838 800
rect 448794 0 448850 800
rect 449806 0 449862 800
rect 450818 0 450874 800
rect 451830 0 451886 800
rect 452842 0 452898 800
rect 453854 0 453910 800
rect 454866 0 454922 800
rect 455878 0 455934 800
rect 456890 0 456946 800
rect 457902 0 457958 800
rect 458914 0 458970 800
rect 459926 0 459982 800
rect 460938 0 460994 800
rect 461950 0 462006 800
rect 462962 0 463018 800
rect 463974 0 464030 800
rect 464986 0 465042 800
rect 465998 0 466054 800
rect 467010 0 467066 800
rect 468022 0 468078 800
rect 469034 0 469090 800
rect 470046 0 470102 800
rect 471058 0 471114 800
rect 472070 0 472126 800
rect 473082 0 473138 800
rect 474094 0 474150 800
rect 475106 0 475162 800
rect 476118 0 476174 800
rect 477130 0 477186 800
rect 478142 0 478198 800
rect 479154 0 479210 800
rect 480166 0 480222 800
rect 481178 0 481234 800
rect 482190 0 482246 800
rect 483202 0 483258 800
rect 484214 0 484270 800
rect 485226 0 485282 800
rect 486238 0 486294 800
rect 487250 0 487306 800
rect 488262 0 488318 800
rect 489274 0 489330 800
rect 490286 0 490342 800
rect 491298 0 491354 800
rect 492310 0 492366 800
rect 493322 0 493378 800
rect 494334 0 494390 800
rect 495346 0 495402 800
rect 496358 0 496414 800
rect 497370 0 497426 800
<< obsm2 >>
rect 938 856 499082 297605
rect 938 70 2446 856
rect 2614 70 3458 856
rect 3626 70 4470 856
rect 4638 70 5482 856
rect 5650 70 6494 856
rect 6662 70 7506 856
rect 7674 70 8518 856
rect 8686 70 9530 856
rect 9698 70 10542 856
rect 10710 70 11554 856
rect 11722 70 12566 856
rect 12734 70 13578 856
rect 13746 70 14590 856
rect 14758 70 15602 856
rect 15770 70 16614 856
rect 16782 70 17626 856
rect 17794 70 18638 856
rect 18806 70 19650 856
rect 19818 70 20662 856
rect 20830 70 21674 856
rect 21842 70 22686 856
rect 22854 70 23698 856
rect 23866 70 24710 856
rect 24878 70 25722 856
rect 25890 70 26734 856
rect 26902 70 27746 856
rect 27914 70 28758 856
rect 28926 70 29770 856
rect 29938 70 30782 856
rect 30950 70 31794 856
rect 31962 70 32806 856
rect 32974 70 33818 856
rect 33986 70 34830 856
rect 34998 70 35842 856
rect 36010 70 36854 856
rect 37022 70 37866 856
rect 38034 70 38878 856
rect 39046 70 39890 856
rect 40058 70 40902 856
rect 41070 70 41914 856
rect 42082 70 42926 856
rect 43094 70 43938 856
rect 44106 70 44950 856
rect 45118 70 45962 856
rect 46130 70 46974 856
rect 47142 70 47986 856
rect 48154 70 48998 856
rect 49166 70 50010 856
rect 50178 70 51022 856
rect 51190 70 52034 856
rect 52202 70 53046 856
rect 53214 70 54058 856
rect 54226 70 55070 856
rect 55238 70 56082 856
rect 56250 70 57094 856
rect 57262 70 58106 856
rect 58274 70 59118 856
rect 59286 70 60130 856
rect 60298 70 61142 856
rect 61310 70 62154 856
rect 62322 70 63166 856
rect 63334 70 64178 856
rect 64346 70 65190 856
rect 65358 70 66202 856
rect 66370 70 67214 856
rect 67382 70 68226 856
rect 68394 70 69238 856
rect 69406 70 70250 856
rect 70418 70 71262 856
rect 71430 70 72274 856
rect 72442 70 73286 856
rect 73454 70 74298 856
rect 74466 70 75310 856
rect 75478 70 76322 856
rect 76490 70 77334 856
rect 77502 70 78346 856
rect 78514 70 79358 856
rect 79526 70 80370 856
rect 80538 70 81382 856
rect 81550 70 82394 856
rect 82562 70 83406 856
rect 83574 70 84418 856
rect 84586 70 85430 856
rect 85598 70 86442 856
rect 86610 70 87454 856
rect 87622 70 88466 856
rect 88634 70 89478 856
rect 89646 70 90490 856
rect 90658 70 91502 856
rect 91670 70 92514 856
rect 92682 70 93526 856
rect 93694 70 94538 856
rect 94706 70 95550 856
rect 95718 70 96562 856
rect 96730 70 97574 856
rect 97742 70 98586 856
rect 98754 70 99598 856
rect 99766 70 100610 856
rect 100778 70 101622 856
rect 101790 70 102634 856
rect 102802 70 103646 856
rect 103814 70 104658 856
rect 104826 70 105670 856
rect 105838 70 106682 856
rect 106850 70 107694 856
rect 107862 70 108706 856
rect 108874 70 109718 856
rect 109886 70 110730 856
rect 110898 70 111742 856
rect 111910 70 112754 856
rect 112922 70 113766 856
rect 113934 70 114778 856
rect 114946 70 115790 856
rect 115958 70 116802 856
rect 116970 70 117814 856
rect 117982 70 118826 856
rect 118994 70 119838 856
rect 120006 70 120850 856
rect 121018 70 121862 856
rect 122030 70 122874 856
rect 123042 70 123886 856
rect 124054 70 124898 856
rect 125066 70 125910 856
rect 126078 70 126922 856
rect 127090 70 127934 856
rect 128102 70 128946 856
rect 129114 70 129958 856
rect 130126 70 130970 856
rect 131138 70 131982 856
rect 132150 70 132994 856
rect 133162 70 134006 856
rect 134174 70 135018 856
rect 135186 70 136030 856
rect 136198 70 137042 856
rect 137210 70 138054 856
rect 138222 70 139066 856
rect 139234 70 140078 856
rect 140246 70 141090 856
rect 141258 70 142102 856
rect 142270 70 143114 856
rect 143282 70 144126 856
rect 144294 70 145138 856
rect 145306 70 146150 856
rect 146318 70 147162 856
rect 147330 70 148174 856
rect 148342 70 149186 856
rect 149354 70 150198 856
rect 150366 70 151210 856
rect 151378 70 152222 856
rect 152390 70 153234 856
rect 153402 70 154246 856
rect 154414 70 155258 856
rect 155426 70 156270 856
rect 156438 70 157282 856
rect 157450 70 158294 856
rect 158462 70 159306 856
rect 159474 70 160318 856
rect 160486 70 161330 856
rect 161498 70 162342 856
rect 162510 70 163354 856
rect 163522 70 164366 856
rect 164534 70 165378 856
rect 165546 70 166390 856
rect 166558 70 167402 856
rect 167570 70 168414 856
rect 168582 70 169426 856
rect 169594 70 170438 856
rect 170606 70 171450 856
rect 171618 70 172462 856
rect 172630 70 173474 856
rect 173642 70 174486 856
rect 174654 70 175498 856
rect 175666 70 176510 856
rect 176678 70 177522 856
rect 177690 70 178534 856
rect 178702 70 179546 856
rect 179714 70 180558 856
rect 180726 70 181570 856
rect 181738 70 182582 856
rect 182750 70 183594 856
rect 183762 70 184606 856
rect 184774 70 185618 856
rect 185786 70 186630 856
rect 186798 70 187642 856
rect 187810 70 188654 856
rect 188822 70 189666 856
rect 189834 70 190678 856
rect 190846 70 191690 856
rect 191858 70 192702 856
rect 192870 70 193714 856
rect 193882 70 194726 856
rect 194894 70 195738 856
rect 195906 70 196750 856
rect 196918 70 197762 856
rect 197930 70 198774 856
rect 198942 70 199786 856
rect 199954 70 200798 856
rect 200966 70 201810 856
rect 201978 70 202822 856
rect 202990 70 203834 856
rect 204002 70 204846 856
rect 205014 70 205858 856
rect 206026 70 206870 856
rect 207038 70 207882 856
rect 208050 70 208894 856
rect 209062 70 209906 856
rect 210074 70 210918 856
rect 211086 70 211930 856
rect 212098 70 212942 856
rect 213110 70 213954 856
rect 214122 70 214966 856
rect 215134 70 215978 856
rect 216146 70 216990 856
rect 217158 70 218002 856
rect 218170 70 219014 856
rect 219182 70 220026 856
rect 220194 70 221038 856
rect 221206 70 222050 856
rect 222218 70 223062 856
rect 223230 70 224074 856
rect 224242 70 225086 856
rect 225254 70 226098 856
rect 226266 70 227110 856
rect 227278 70 228122 856
rect 228290 70 229134 856
rect 229302 70 230146 856
rect 230314 70 231158 856
rect 231326 70 232170 856
rect 232338 70 233182 856
rect 233350 70 234194 856
rect 234362 70 235206 856
rect 235374 70 236218 856
rect 236386 70 237230 856
rect 237398 70 238242 856
rect 238410 70 239254 856
rect 239422 70 240266 856
rect 240434 70 241278 856
rect 241446 70 242290 856
rect 242458 70 243302 856
rect 243470 70 244314 856
rect 244482 70 245326 856
rect 245494 70 246338 856
rect 246506 70 247350 856
rect 247518 70 248362 856
rect 248530 70 249374 856
rect 249542 70 250386 856
rect 250554 70 251398 856
rect 251566 70 252410 856
rect 252578 70 253422 856
rect 253590 70 254434 856
rect 254602 70 255446 856
rect 255614 70 256458 856
rect 256626 70 257470 856
rect 257638 70 258482 856
rect 258650 70 259494 856
rect 259662 70 260506 856
rect 260674 70 261518 856
rect 261686 70 262530 856
rect 262698 70 263542 856
rect 263710 70 264554 856
rect 264722 70 265566 856
rect 265734 70 266578 856
rect 266746 70 267590 856
rect 267758 70 268602 856
rect 268770 70 269614 856
rect 269782 70 270626 856
rect 270794 70 271638 856
rect 271806 70 272650 856
rect 272818 70 273662 856
rect 273830 70 274674 856
rect 274842 70 275686 856
rect 275854 70 276698 856
rect 276866 70 277710 856
rect 277878 70 278722 856
rect 278890 70 279734 856
rect 279902 70 280746 856
rect 280914 70 281758 856
rect 281926 70 282770 856
rect 282938 70 283782 856
rect 283950 70 284794 856
rect 284962 70 285806 856
rect 285974 70 286818 856
rect 286986 70 287830 856
rect 287998 70 288842 856
rect 289010 70 289854 856
rect 290022 70 290866 856
rect 291034 70 291878 856
rect 292046 70 292890 856
rect 293058 70 293902 856
rect 294070 70 294914 856
rect 295082 70 295926 856
rect 296094 70 296938 856
rect 297106 70 297950 856
rect 298118 70 298962 856
rect 299130 70 299974 856
rect 300142 70 300986 856
rect 301154 70 301998 856
rect 302166 70 303010 856
rect 303178 70 304022 856
rect 304190 70 305034 856
rect 305202 70 306046 856
rect 306214 70 307058 856
rect 307226 70 308070 856
rect 308238 70 309082 856
rect 309250 70 310094 856
rect 310262 70 311106 856
rect 311274 70 312118 856
rect 312286 70 313130 856
rect 313298 70 314142 856
rect 314310 70 315154 856
rect 315322 70 316166 856
rect 316334 70 317178 856
rect 317346 70 318190 856
rect 318358 70 319202 856
rect 319370 70 320214 856
rect 320382 70 321226 856
rect 321394 70 322238 856
rect 322406 70 323250 856
rect 323418 70 324262 856
rect 324430 70 325274 856
rect 325442 70 326286 856
rect 326454 70 327298 856
rect 327466 70 328310 856
rect 328478 70 329322 856
rect 329490 70 330334 856
rect 330502 70 331346 856
rect 331514 70 332358 856
rect 332526 70 333370 856
rect 333538 70 334382 856
rect 334550 70 335394 856
rect 335562 70 336406 856
rect 336574 70 337418 856
rect 337586 70 338430 856
rect 338598 70 339442 856
rect 339610 70 340454 856
rect 340622 70 341466 856
rect 341634 70 342478 856
rect 342646 70 343490 856
rect 343658 70 344502 856
rect 344670 70 345514 856
rect 345682 70 346526 856
rect 346694 70 347538 856
rect 347706 70 348550 856
rect 348718 70 349562 856
rect 349730 70 350574 856
rect 350742 70 351586 856
rect 351754 70 352598 856
rect 352766 70 353610 856
rect 353778 70 354622 856
rect 354790 70 355634 856
rect 355802 70 356646 856
rect 356814 70 357658 856
rect 357826 70 358670 856
rect 358838 70 359682 856
rect 359850 70 360694 856
rect 360862 70 361706 856
rect 361874 70 362718 856
rect 362886 70 363730 856
rect 363898 70 364742 856
rect 364910 70 365754 856
rect 365922 70 366766 856
rect 366934 70 367778 856
rect 367946 70 368790 856
rect 368958 70 369802 856
rect 369970 70 370814 856
rect 370982 70 371826 856
rect 371994 70 372838 856
rect 373006 70 373850 856
rect 374018 70 374862 856
rect 375030 70 375874 856
rect 376042 70 376886 856
rect 377054 70 377898 856
rect 378066 70 378910 856
rect 379078 70 379922 856
rect 380090 70 380934 856
rect 381102 70 381946 856
rect 382114 70 382958 856
rect 383126 70 383970 856
rect 384138 70 384982 856
rect 385150 70 385994 856
rect 386162 70 387006 856
rect 387174 70 388018 856
rect 388186 70 389030 856
rect 389198 70 390042 856
rect 390210 70 391054 856
rect 391222 70 392066 856
rect 392234 70 393078 856
rect 393246 70 394090 856
rect 394258 70 395102 856
rect 395270 70 396114 856
rect 396282 70 397126 856
rect 397294 70 398138 856
rect 398306 70 399150 856
rect 399318 70 400162 856
rect 400330 70 401174 856
rect 401342 70 402186 856
rect 402354 70 403198 856
rect 403366 70 404210 856
rect 404378 70 405222 856
rect 405390 70 406234 856
rect 406402 70 407246 856
rect 407414 70 408258 856
rect 408426 70 409270 856
rect 409438 70 410282 856
rect 410450 70 411294 856
rect 411462 70 412306 856
rect 412474 70 413318 856
rect 413486 70 414330 856
rect 414498 70 415342 856
rect 415510 70 416354 856
rect 416522 70 417366 856
rect 417534 70 418378 856
rect 418546 70 419390 856
rect 419558 70 420402 856
rect 420570 70 421414 856
rect 421582 70 422426 856
rect 422594 70 423438 856
rect 423606 70 424450 856
rect 424618 70 425462 856
rect 425630 70 426474 856
rect 426642 70 427486 856
rect 427654 70 428498 856
rect 428666 70 429510 856
rect 429678 70 430522 856
rect 430690 70 431534 856
rect 431702 70 432546 856
rect 432714 70 433558 856
rect 433726 70 434570 856
rect 434738 70 435582 856
rect 435750 70 436594 856
rect 436762 70 437606 856
rect 437774 70 438618 856
rect 438786 70 439630 856
rect 439798 70 440642 856
rect 440810 70 441654 856
rect 441822 70 442666 856
rect 442834 70 443678 856
rect 443846 70 444690 856
rect 444858 70 445702 856
rect 445870 70 446714 856
rect 446882 70 447726 856
rect 447894 70 448738 856
rect 448906 70 449750 856
rect 449918 70 450762 856
rect 450930 70 451774 856
rect 451942 70 452786 856
rect 452954 70 453798 856
rect 453966 70 454810 856
rect 454978 70 455822 856
rect 455990 70 456834 856
rect 457002 70 457846 856
rect 458014 70 458858 856
rect 459026 70 459870 856
rect 460038 70 460882 856
rect 461050 70 461894 856
rect 462062 70 462906 856
rect 463074 70 463918 856
rect 464086 70 464930 856
rect 465098 70 465942 856
rect 466110 70 466954 856
rect 467122 70 467966 856
rect 468134 70 468978 856
rect 469146 70 469990 856
rect 470158 70 471002 856
rect 471170 70 472014 856
rect 472182 70 473026 856
rect 473194 70 474038 856
rect 474206 70 475050 856
rect 475218 70 476062 856
rect 476230 70 477074 856
rect 477242 70 478086 856
rect 478254 70 479098 856
rect 479266 70 480110 856
rect 480278 70 481122 856
rect 481290 70 482134 856
rect 482302 70 483146 856
rect 483314 70 484158 856
rect 484326 70 485170 856
rect 485338 70 486182 856
rect 486350 70 487194 856
rect 487362 70 488206 856
rect 488374 70 489218 856
rect 489386 70 490230 856
rect 490398 70 491242 856
rect 491410 70 492254 856
rect 492422 70 493266 856
rect 493434 70 494278 856
rect 494446 70 495290 856
rect 495458 70 496302 856
rect 496470 70 497314 856
rect 497482 70 499082 856
<< metal3 >>
rect 0 292272 800 292392
rect 499200 292272 500000 292392
rect 0 279896 800 280016
rect 499200 279896 500000 280016
rect 0 267520 800 267640
rect 499200 267520 500000 267640
rect 0 255144 800 255264
rect 499200 255144 500000 255264
rect 0 242768 800 242888
rect 499200 242768 500000 242888
rect 0 230392 800 230512
rect 499200 230392 500000 230512
rect 0 218016 800 218136
rect 499200 218016 500000 218136
rect 0 205640 800 205760
rect 499200 205640 500000 205760
rect 0 193264 800 193384
rect 499200 193264 500000 193384
rect 0 180888 800 181008
rect 499200 180888 500000 181008
rect 0 168512 800 168632
rect 499200 168512 500000 168632
rect 0 156136 800 156256
rect 499200 156136 500000 156256
rect 0 143760 800 143880
rect 499200 143760 500000 143880
rect 0 131384 800 131504
rect 499200 131384 500000 131504
rect 0 119008 800 119128
rect 499200 119008 500000 119128
rect 0 106632 800 106752
rect 499200 106632 500000 106752
rect 0 94256 800 94376
rect 499200 94256 500000 94376
rect 0 81880 800 82000
rect 499200 81880 500000 82000
rect 0 69504 800 69624
rect 499200 69504 500000 69624
rect 0 57128 800 57248
rect 499200 57128 500000 57248
rect 0 44752 800 44872
rect 499200 44752 500000 44872
rect 0 32376 800 32496
rect 499200 32376 500000 32496
rect 0 20000 800 20120
rect 499200 20000 500000 20120
rect 0 7624 800 7744
rect 499200 7624 500000 7744
<< obsm3 >>
rect 800 292472 499200 297601
rect 880 292192 499120 292472
rect 800 280096 499200 292192
rect 880 279816 499120 280096
rect 800 267720 499200 279816
rect 880 267440 499120 267720
rect 800 255344 499200 267440
rect 880 255064 499120 255344
rect 800 242968 499200 255064
rect 880 242688 499120 242968
rect 800 230592 499200 242688
rect 880 230312 499120 230592
rect 800 218216 499200 230312
rect 880 217936 499120 218216
rect 800 205840 499200 217936
rect 880 205560 499120 205840
rect 800 193464 499200 205560
rect 880 193184 499120 193464
rect 800 181088 499200 193184
rect 880 180808 499120 181088
rect 800 168712 499200 180808
rect 880 168432 499120 168712
rect 800 156336 499200 168432
rect 880 156056 499120 156336
rect 800 143960 499200 156056
rect 880 143680 499120 143960
rect 800 131584 499200 143680
rect 880 131304 499120 131584
rect 800 119208 499200 131304
rect 880 118928 499120 119208
rect 800 106832 499200 118928
rect 880 106552 499120 106832
rect 800 94456 499200 106552
rect 880 94176 499120 94456
rect 800 82080 499200 94176
rect 880 81800 499120 82080
rect 800 69704 499200 81800
rect 880 69424 499120 69704
rect 800 57328 499200 69424
rect 880 57048 499120 57328
rect 800 44952 499200 57048
rect 880 44672 499120 44952
rect 800 32576 499200 44672
rect 880 32296 499120 32576
rect 800 20200 499200 32296
rect 880 19920 499120 20200
rect 800 7824 499200 19920
rect 880 7544 499120 7824
rect 800 2143 499200 7544
<< metal4 >>
rect 4208 2128 4528 297616
rect 19568 2128 19888 297616
rect 34928 2128 35248 297616
rect 50288 2128 50608 297616
rect 65648 2128 65968 297616
rect 81008 2128 81328 297616
rect 96368 2128 96688 297616
rect 111728 2128 112048 297616
rect 127088 2128 127408 297616
rect 142448 2128 142768 297616
rect 157808 2128 158128 297616
rect 173168 2128 173488 297616
rect 188528 2128 188848 297616
rect 203888 2128 204208 297616
rect 219248 2128 219568 297616
rect 234608 2128 234928 297616
rect 249968 2128 250288 297616
rect 265328 2128 265648 297616
rect 280688 2128 281008 297616
rect 296048 2128 296368 297616
rect 311408 2128 311728 297616
rect 326768 2128 327088 297616
rect 342128 2128 342448 297616
rect 357488 2128 357808 297616
rect 372848 2128 373168 297616
rect 388208 2128 388528 297616
rect 403568 2128 403888 297616
rect 418928 2128 419248 297616
rect 434288 2128 434608 297616
rect 449648 2128 449968 297616
rect 465008 2128 465328 297616
rect 480368 2128 480688 297616
rect 495728 2128 496048 297616
<< labels >>
rlabel metal3 s 499200 7624 500000 7744 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 0 218016 800 218136 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 0 180888 800 181008 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 0 143760 800 143880 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 0 106632 800 106752 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 0 69504 800 69624 6 io_in[14]
port 6 nsew signal input
rlabel metal3 s 0 32376 800 32496 6 io_in[15]
port 7 nsew signal input
rlabel metal3 s 499200 44752 500000 44872 6 io_in[1]
port 8 nsew signal input
rlabel metal3 s 499200 81880 500000 82000 6 io_in[2]
port 9 nsew signal input
rlabel metal3 s 499200 119008 500000 119128 6 io_in[3]
port 10 nsew signal input
rlabel metal3 s 499200 156136 500000 156256 6 io_in[4]
port 11 nsew signal input
rlabel metal3 s 499200 193264 500000 193384 6 io_in[5]
port 12 nsew signal input
rlabel metal3 s 499200 230392 500000 230512 6 io_in[6]
port 13 nsew signal input
rlabel metal3 s 499200 267520 500000 267640 6 io_in[7]
port 14 nsew signal input
rlabel metal3 s 0 292272 800 292392 6 io_in[8]
port 15 nsew signal input
rlabel metal3 s 0 255144 800 255264 6 io_in[9]
port 16 nsew signal input
rlabel metal3 s 499200 32376 500000 32496 6 io_oeb[0]
port 17 nsew signal output
rlabel metal3 s 0 193264 800 193384 6 io_oeb[10]
port 18 nsew signal output
rlabel metal3 s 0 156136 800 156256 6 io_oeb[11]
port 19 nsew signal output
rlabel metal3 s 0 119008 800 119128 6 io_oeb[12]
port 20 nsew signal output
rlabel metal3 s 0 81880 800 82000 6 io_oeb[13]
port 21 nsew signal output
rlabel metal3 s 0 44752 800 44872 6 io_oeb[14]
port 22 nsew signal output
rlabel metal3 s 0 7624 800 7744 6 io_oeb[15]
port 23 nsew signal output
rlabel metal3 s 499200 69504 500000 69624 6 io_oeb[1]
port 24 nsew signal output
rlabel metal3 s 499200 106632 500000 106752 6 io_oeb[2]
port 25 nsew signal output
rlabel metal3 s 499200 143760 500000 143880 6 io_oeb[3]
port 26 nsew signal output
rlabel metal3 s 499200 180888 500000 181008 6 io_oeb[4]
port 27 nsew signal output
rlabel metal3 s 499200 218016 500000 218136 6 io_oeb[5]
port 28 nsew signal output
rlabel metal3 s 499200 255144 500000 255264 6 io_oeb[6]
port 29 nsew signal output
rlabel metal3 s 499200 292272 500000 292392 6 io_oeb[7]
port 30 nsew signal output
rlabel metal3 s 0 267520 800 267640 6 io_oeb[8]
port 31 nsew signal output
rlabel metal3 s 0 230392 800 230512 6 io_oeb[9]
port 32 nsew signal output
rlabel metal3 s 499200 20000 500000 20120 6 io_out[0]
port 33 nsew signal output
rlabel metal3 s 0 205640 800 205760 6 io_out[10]
port 34 nsew signal output
rlabel metal3 s 0 168512 800 168632 6 io_out[11]
port 35 nsew signal output
rlabel metal3 s 0 131384 800 131504 6 io_out[12]
port 36 nsew signal output
rlabel metal3 s 0 94256 800 94376 6 io_out[13]
port 37 nsew signal output
rlabel metal3 s 0 57128 800 57248 6 io_out[14]
port 38 nsew signal output
rlabel metal3 s 0 20000 800 20120 6 io_out[15]
port 39 nsew signal output
rlabel metal3 s 499200 57128 500000 57248 6 io_out[1]
port 40 nsew signal output
rlabel metal3 s 499200 94256 500000 94376 6 io_out[2]
port 41 nsew signal output
rlabel metal3 s 499200 131384 500000 131504 6 io_out[3]
port 42 nsew signal output
rlabel metal3 s 499200 168512 500000 168632 6 io_out[4]
port 43 nsew signal output
rlabel metal3 s 499200 205640 500000 205760 6 io_out[5]
port 44 nsew signal output
rlabel metal3 s 499200 242768 500000 242888 6 io_out[6]
port 45 nsew signal output
rlabel metal3 s 499200 279896 500000 280016 6 io_out[7]
port 46 nsew signal output
rlabel metal3 s 0 279896 800 280016 6 io_out[8]
port 47 nsew signal output
rlabel metal3 s 0 242768 800 242888 6 io_out[9]
port 48 nsew signal output
rlabel metal2 s 109774 0 109830 800 6 la_data_in[0]
port 49 nsew signal input
rlabel metal2 s 413374 0 413430 800 6 la_data_in[100]
port 50 nsew signal input
rlabel metal2 s 416410 0 416466 800 6 la_data_in[101]
port 51 nsew signal input
rlabel metal2 s 419446 0 419502 800 6 la_data_in[102]
port 52 nsew signal input
rlabel metal2 s 422482 0 422538 800 6 la_data_in[103]
port 53 nsew signal input
rlabel metal2 s 425518 0 425574 800 6 la_data_in[104]
port 54 nsew signal input
rlabel metal2 s 428554 0 428610 800 6 la_data_in[105]
port 55 nsew signal input
rlabel metal2 s 431590 0 431646 800 6 la_data_in[106]
port 56 nsew signal input
rlabel metal2 s 434626 0 434682 800 6 la_data_in[107]
port 57 nsew signal input
rlabel metal2 s 437662 0 437718 800 6 la_data_in[108]
port 58 nsew signal input
rlabel metal2 s 440698 0 440754 800 6 la_data_in[109]
port 59 nsew signal input
rlabel metal2 s 140134 0 140190 800 6 la_data_in[10]
port 60 nsew signal input
rlabel metal2 s 443734 0 443790 800 6 la_data_in[110]
port 61 nsew signal input
rlabel metal2 s 446770 0 446826 800 6 la_data_in[111]
port 62 nsew signal input
rlabel metal2 s 449806 0 449862 800 6 la_data_in[112]
port 63 nsew signal input
rlabel metal2 s 452842 0 452898 800 6 la_data_in[113]
port 64 nsew signal input
rlabel metal2 s 455878 0 455934 800 6 la_data_in[114]
port 65 nsew signal input
rlabel metal2 s 458914 0 458970 800 6 la_data_in[115]
port 66 nsew signal input
rlabel metal2 s 461950 0 462006 800 6 la_data_in[116]
port 67 nsew signal input
rlabel metal2 s 464986 0 465042 800 6 la_data_in[117]
port 68 nsew signal input
rlabel metal2 s 468022 0 468078 800 6 la_data_in[118]
port 69 nsew signal input
rlabel metal2 s 471058 0 471114 800 6 la_data_in[119]
port 70 nsew signal input
rlabel metal2 s 143170 0 143226 800 6 la_data_in[11]
port 71 nsew signal input
rlabel metal2 s 474094 0 474150 800 6 la_data_in[120]
port 72 nsew signal input
rlabel metal2 s 477130 0 477186 800 6 la_data_in[121]
port 73 nsew signal input
rlabel metal2 s 480166 0 480222 800 6 la_data_in[122]
port 74 nsew signal input
rlabel metal2 s 483202 0 483258 800 6 la_data_in[123]
port 75 nsew signal input
rlabel metal2 s 486238 0 486294 800 6 la_data_in[124]
port 76 nsew signal input
rlabel metal2 s 489274 0 489330 800 6 la_data_in[125]
port 77 nsew signal input
rlabel metal2 s 492310 0 492366 800 6 la_data_in[126]
port 78 nsew signal input
rlabel metal2 s 495346 0 495402 800 6 la_data_in[127]
port 79 nsew signal input
rlabel metal2 s 146206 0 146262 800 6 la_data_in[12]
port 80 nsew signal input
rlabel metal2 s 149242 0 149298 800 6 la_data_in[13]
port 81 nsew signal input
rlabel metal2 s 152278 0 152334 800 6 la_data_in[14]
port 82 nsew signal input
rlabel metal2 s 155314 0 155370 800 6 la_data_in[15]
port 83 nsew signal input
rlabel metal2 s 158350 0 158406 800 6 la_data_in[16]
port 84 nsew signal input
rlabel metal2 s 161386 0 161442 800 6 la_data_in[17]
port 85 nsew signal input
rlabel metal2 s 164422 0 164478 800 6 la_data_in[18]
port 86 nsew signal input
rlabel metal2 s 167458 0 167514 800 6 la_data_in[19]
port 87 nsew signal input
rlabel metal2 s 112810 0 112866 800 6 la_data_in[1]
port 88 nsew signal input
rlabel metal2 s 170494 0 170550 800 6 la_data_in[20]
port 89 nsew signal input
rlabel metal2 s 173530 0 173586 800 6 la_data_in[21]
port 90 nsew signal input
rlabel metal2 s 176566 0 176622 800 6 la_data_in[22]
port 91 nsew signal input
rlabel metal2 s 179602 0 179658 800 6 la_data_in[23]
port 92 nsew signal input
rlabel metal2 s 182638 0 182694 800 6 la_data_in[24]
port 93 nsew signal input
rlabel metal2 s 185674 0 185730 800 6 la_data_in[25]
port 94 nsew signal input
rlabel metal2 s 188710 0 188766 800 6 la_data_in[26]
port 95 nsew signal input
rlabel metal2 s 191746 0 191802 800 6 la_data_in[27]
port 96 nsew signal input
rlabel metal2 s 194782 0 194838 800 6 la_data_in[28]
port 97 nsew signal input
rlabel metal2 s 197818 0 197874 800 6 la_data_in[29]
port 98 nsew signal input
rlabel metal2 s 115846 0 115902 800 6 la_data_in[2]
port 99 nsew signal input
rlabel metal2 s 200854 0 200910 800 6 la_data_in[30]
port 100 nsew signal input
rlabel metal2 s 203890 0 203946 800 6 la_data_in[31]
port 101 nsew signal input
rlabel metal2 s 206926 0 206982 800 6 la_data_in[32]
port 102 nsew signal input
rlabel metal2 s 209962 0 210018 800 6 la_data_in[33]
port 103 nsew signal input
rlabel metal2 s 212998 0 213054 800 6 la_data_in[34]
port 104 nsew signal input
rlabel metal2 s 216034 0 216090 800 6 la_data_in[35]
port 105 nsew signal input
rlabel metal2 s 219070 0 219126 800 6 la_data_in[36]
port 106 nsew signal input
rlabel metal2 s 222106 0 222162 800 6 la_data_in[37]
port 107 nsew signal input
rlabel metal2 s 225142 0 225198 800 6 la_data_in[38]
port 108 nsew signal input
rlabel metal2 s 228178 0 228234 800 6 la_data_in[39]
port 109 nsew signal input
rlabel metal2 s 118882 0 118938 800 6 la_data_in[3]
port 110 nsew signal input
rlabel metal2 s 231214 0 231270 800 6 la_data_in[40]
port 111 nsew signal input
rlabel metal2 s 234250 0 234306 800 6 la_data_in[41]
port 112 nsew signal input
rlabel metal2 s 237286 0 237342 800 6 la_data_in[42]
port 113 nsew signal input
rlabel metal2 s 240322 0 240378 800 6 la_data_in[43]
port 114 nsew signal input
rlabel metal2 s 243358 0 243414 800 6 la_data_in[44]
port 115 nsew signal input
rlabel metal2 s 246394 0 246450 800 6 la_data_in[45]
port 116 nsew signal input
rlabel metal2 s 249430 0 249486 800 6 la_data_in[46]
port 117 nsew signal input
rlabel metal2 s 252466 0 252522 800 6 la_data_in[47]
port 118 nsew signal input
rlabel metal2 s 255502 0 255558 800 6 la_data_in[48]
port 119 nsew signal input
rlabel metal2 s 258538 0 258594 800 6 la_data_in[49]
port 120 nsew signal input
rlabel metal2 s 121918 0 121974 800 6 la_data_in[4]
port 121 nsew signal input
rlabel metal2 s 261574 0 261630 800 6 la_data_in[50]
port 122 nsew signal input
rlabel metal2 s 264610 0 264666 800 6 la_data_in[51]
port 123 nsew signal input
rlabel metal2 s 267646 0 267702 800 6 la_data_in[52]
port 124 nsew signal input
rlabel metal2 s 270682 0 270738 800 6 la_data_in[53]
port 125 nsew signal input
rlabel metal2 s 273718 0 273774 800 6 la_data_in[54]
port 126 nsew signal input
rlabel metal2 s 276754 0 276810 800 6 la_data_in[55]
port 127 nsew signal input
rlabel metal2 s 279790 0 279846 800 6 la_data_in[56]
port 128 nsew signal input
rlabel metal2 s 282826 0 282882 800 6 la_data_in[57]
port 129 nsew signal input
rlabel metal2 s 285862 0 285918 800 6 la_data_in[58]
port 130 nsew signal input
rlabel metal2 s 288898 0 288954 800 6 la_data_in[59]
port 131 nsew signal input
rlabel metal2 s 124954 0 125010 800 6 la_data_in[5]
port 132 nsew signal input
rlabel metal2 s 291934 0 291990 800 6 la_data_in[60]
port 133 nsew signal input
rlabel metal2 s 294970 0 295026 800 6 la_data_in[61]
port 134 nsew signal input
rlabel metal2 s 298006 0 298062 800 6 la_data_in[62]
port 135 nsew signal input
rlabel metal2 s 301042 0 301098 800 6 la_data_in[63]
port 136 nsew signal input
rlabel metal2 s 304078 0 304134 800 6 la_data_in[64]
port 137 nsew signal input
rlabel metal2 s 307114 0 307170 800 6 la_data_in[65]
port 138 nsew signal input
rlabel metal2 s 310150 0 310206 800 6 la_data_in[66]
port 139 nsew signal input
rlabel metal2 s 313186 0 313242 800 6 la_data_in[67]
port 140 nsew signal input
rlabel metal2 s 316222 0 316278 800 6 la_data_in[68]
port 141 nsew signal input
rlabel metal2 s 319258 0 319314 800 6 la_data_in[69]
port 142 nsew signal input
rlabel metal2 s 127990 0 128046 800 6 la_data_in[6]
port 143 nsew signal input
rlabel metal2 s 322294 0 322350 800 6 la_data_in[70]
port 144 nsew signal input
rlabel metal2 s 325330 0 325386 800 6 la_data_in[71]
port 145 nsew signal input
rlabel metal2 s 328366 0 328422 800 6 la_data_in[72]
port 146 nsew signal input
rlabel metal2 s 331402 0 331458 800 6 la_data_in[73]
port 147 nsew signal input
rlabel metal2 s 334438 0 334494 800 6 la_data_in[74]
port 148 nsew signal input
rlabel metal2 s 337474 0 337530 800 6 la_data_in[75]
port 149 nsew signal input
rlabel metal2 s 340510 0 340566 800 6 la_data_in[76]
port 150 nsew signal input
rlabel metal2 s 343546 0 343602 800 6 la_data_in[77]
port 151 nsew signal input
rlabel metal2 s 346582 0 346638 800 6 la_data_in[78]
port 152 nsew signal input
rlabel metal2 s 349618 0 349674 800 6 la_data_in[79]
port 153 nsew signal input
rlabel metal2 s 131026 0 131082 800 6 la_data_in[7]
port 154 nsew signal input
rlabel metal2 s 352654 0 352710 800 6 la_data_in[80]
port 155 nsew signal input
rlabel metal2 s 355690 0 355746 800 6 la_data_in[81]
port 156 nsew signal input
rlabel metal2 s 358726 0 358782 800 6 la_data_in[82]
port 157 nsew signal input
rlabel metal2 s 361762 0 361818 800 6 la_data_in[83]
port 158 nsew signal input
rlabel metal2 s 364798 0 364854 800 6 la_data_in[84]
port 159 nsew signal input
rlabel metal2 s 367834 0 367890 800 6 la_data_in[85]
port 160 nsew signal input
rlabel metal2 s 370870 0 370926 800 6 la_data_in[86]
port 161 nsew signal input
rlabel metal2 s 373906 0 373962 800 6 la_data_in[87]
port 162 nsew signal input
rlabel metal2 s 376942 0 376998 800 6 la_data_in[88]
port 163 nsew signal input
rlabel metal2 s 379978 0 380034 800 6 la_data_in[89]
port 164 nsew signal input
rlabel metal2 s 134062 0 134118 800 6 la_data_in[8]
port 165 nsew signal input
rlabel metal2 s 383014 0 383070 800 6 la_data_in[90]
port 166 nsew signal input
rlabel metal2 s 386050 0 386106 800 6 la_data_in[91]
port 167 nsew signal input
rlabel metal2 s 389086 0 389142 800 6 la_data_in[92]
port 168 nsew signal input
rlabel metal2 s 392122 0 392178 800 6 la_data_in[93]
port 169 nsew signal input
rlabel metal2 s 395158 0 395214 800 6 la_data_in[94]
port 170 nsew signal input
rlabel metal2 s 398194 0 398250 800 6 la_data_in[95]
port 171 nsew signal input
rlabel metal2 s 401230 0 401286 800 6 la_data_in[96]
port 172 nsew signal input
rlabel metal2 s 404266 0 404322 800 6 la_data_in[97]
port 173 nsew signal input
rlabel metal2 s 407302 0 407358 800 6 la_data_in[98]
port 174 nsew signal input
rlabel metal2 s 410338 0 410394 800 6 la_data_in[99]
port 175 nsew signal input
rlabel metal2 s 137098 0 137154 800 6 la_data_in[9]
port 176 nsew signal input
rlabel metal2 s 110786 0 110842 800 6 la_data_out[0]
port 177 nsew signal output
rlabel metal2 s 414386 0 414442 800 6 la_data_out[100]
port 178 nsew signal output
rlabel metal2 s 417422 0 417478 800 6 la_data_out[101]
port 179 nsew signal output
rlabel metal2 s 420458 0 420514 800 6 la_data_out[102]
port 180 nsew signal output
rlabel metal2 s 423494 0 423550 800 6 la_data_out[103]
port 181 nsew signal output
rlabel metal2 s 426530 0 426586 800 6 la_data_out[104]
port 182 nsew signal output
rlabel metal2 s 429566 0 429622 800 6 la_data_out[105]
port 183 nsew signal output
rlabel metal2 s 432602 0 432658 800 6 la_data_out[106]
port 184 nsew signal output
rlabel metal2 s 435638 0 435694 800 6 la_data_out[107]
port 185 nsew signal output
rlabel metal2 s 438674 0 438730 800 6 la_data_out[108]
port 186 nsew signal output
rlabel metal2 s 441710 0 441766 800 6 la_data_out[109]
port 187 nsew signal output
rlabel metal2 s 141146 0 141202 800 6 la_data_out[10]
port 188 nsew signal output
rlabel metal2 s 444746 0 444802 800 6 la_data_out[110]
port 189 nsew signal output
rlabel metal2 s 447782 0 447838 800 6 la_data_out[111]
port 190 nsew signal output
rlabel metal2 s 450818 0 450874 800 6 la_data_out[112]
port 191 nsew signal output
rlabel metal2 s 453854 0 453910 800 6 la_data_out[113]
port 192 nsew signal output
rlabel metal2 s 456890 0 456946 800 6 la_data_out[114]
port 193 nsew signal output
rlabel metal2 s 459926 0 459982 800 6 la_data_out[115]
port 194 nsew signal output
rlabel metal2 s 462962 0 463018 800 6 la_data_out[116]
port 195 nsew signal output
rlabel metal2 s 465998 0 466054 800 6 la_data_out[117]
port 196 nsew signal output
rlabel metal2 s 469034 0 469090 800 6 la_data_out[118]
port 197 nsew signal output
rlabel metal2 s 472070 0 472126 800 6 la_data_out[119]
port 198 nsew signal output
rlabel metal2 s 144182 0 144238 800 6 la_data_out[11]
port 199 nsew signal output
rlabel metal2 s 475106 0 475162 800 6 la_data_out[120]
port 200 nsew signal output
rlabel metal2 s 478142 0 478198 800 6 la_data_out[121]
port 201 nsew signal output
rlabel metal2 s 481178 0 481234 800 6 la_data_out[122]
port 202 nsew signal output
rlabel metal2 s 484214 0 484270 800 6 la_data_out[123]
port 203 nsew signal output
rlabel metal2 s 487250 0 487306 800 6 la_data_out[124]
port 204 nsew signal output
rlabel metal2 s 490286 0 490342 800 6 la_data_out[125]
port 205 nsew signal output
rlabel metal2 s 493322 0 493378 800 6 la_data_out[126]
port 206 nsew signal output
rlabel metal2 s 496358 0 496414 800 6 la_data_out[127]
port 207 nsew signal output
rlabel metal2 s 147218 0 147274 800 6 la_data_out[12]
port 208 nsew signal output
rlabel metal2 s 150254 0 150310 800 6 la_data_out[13]
port 209 nsew signal output
rlabel metal2 s 153290 0 153346 800 6 la_data_out[14]
port 210 nsew signal output
rlabel metal2 s 156326 0 156382 800 6 la_data_out[15]
port 211 nsew signal output
rlabel metal2 s 159362 0 159418 800 6 la_data_out[16]
port 212 nsew signal output
rlabel metal2 s 162398 0 162454 800 6 la_data_out[17]
port 213 nsew signal output
rlabel metal2 s 165434 0 165490 800 6 la_data_out[18]
port 214 nsew signal output
rlabel metal2 s 168470 0 168526 800 6 la_data_out[19]
port 215 nsew signal output
rlabel metal2 s 113822 0 113878 800 6 la_data_out[1]
port 216 nsew signal output
rlabel metal2 s 171506 0 171562 800 6 la_data_out[20]
port 217 nsew signal output
rlabel metal2 s 174542 0 174598 800 6 la_data_out[21]
port 218 nsew signal output
rlabel metal2 s 177578 0 177634 800 6 la_data_out[22]
port 219 nsew signal output
rlabel metal2 s 180614 0 180670 800 6 la_data_out[23]
port 220 nsew signal output
rlabel metal2 s 183650 0 183706 800 6 la_data_out[24]
port 221 nsew signal output
rlabel metal2 s 186686 0 186742 800 6 la_data_out[25]
port 222 nsew signal output
rlabel metal2 s 189722 0 189778 800 6 la_data_out[26]
port 223 nsew signal output
rlabel metal2 s 192758 0 192814 800 6 la_data_out[27]
port 224 nsew signal output
rlabel metal2 s 195794 0 195850 800 6 la_data_out[28]
port 225 nsew signal output
rlabel metal2 s 198830 0 198886 800 6 la_data_out[29]
port 226 nsew signal output
rlabel metal2 s 116858 0 116914 800 6 la_data_out[2]
port 227 nsew signal output
rlabel metal2 s 201866 0 201922 800 6 la_data_out[30]
port 228 nsew signal output
rlabel metal2 s 204902 0 204958 800 6 la_data_out[31]
port 229 nsew signal output
rlabel metal2 s 207938 0 207994 800 6 la_data_out[32]
port 230 nsew signal output
rlabel metal2 s 210974 0 211030 800 6 la_data_out[33]
port 231 nsew signal output
rlabel metal2 s 214010 0 214066 800 6 la_data_out[34]
port 232 nsew signal output
rlabel metal2 s 217046 0 217102 800 6 la_data_out[35]
port 233 nsew signal output
rlabel metal2 s 220082 0 220138 800 6 la_data_out[36]
port 234 nsew signal output
rlabel metal2 s 223118 0 223174 800 6 la_data_out[37]
port 235 nsew signal output
rlabel metal2 s 226154 0 226210 800 6 la_data_out[38]
port 236 nsew signal output
rlabel metal2 s 229190 0 229246 800 6 la_data_out[39]
port 237 nsew signal output
rlabel metal2 s 119894 0 119950 800 6 la_data_out[3]
port 238 nsew signal output
rlabel metal2 s 232226 0 232282 800 6 la_data_out[40]
port 239 nsew signal output
rlabel metal2 s 235262 0 235318 800 6 la_data_out[41]
port 240 nsew signal output
rlabel metal2 s 238298 0 238354 800 6 la_data_out[42]
port 241 nsew signal output
rlabel metal2 s 241334 0 241390 800 6 la_data_out[43]
port 242 nsew signal output
rlabel metal2 s 244370 0 244426 800 6 la_data_out[44]
port 243 nsew signal output
rlabel metal2 s 247406 0 247462 800 6 la_data_out[45]
port 244 nsew signal output
rlabel metal2 s 250442 0 250498 800 6 la_data_out[46]
port 245 nsew signal output
rlabel metal2 s 253478 0 253534 800 6 la_data_out[47]
port 246 nsew signal output
rlabel metal2 s 256514 0 256570 800 6 la_data_out[48]
port 247 nsew signal output
rlabel metal2 s 259550 0 259606 800 6 la_data_out[49]
port 248 nsew signal output
rlabel metal2 s 122930 0 122986 800 6 la_data_out[4]
port 249 nsew signal output
rlabel metal2 s 262586 0 262642 800 6 la_data_out[50]
port 250 nsew signal output
rlabel metal2 s 265622 0 265678 800 6 la_data_out[51]
port 251 nsew signal output
rlabel metal2 s 268658 0 268714 800 6 la_data_out[52]
port 252 nsew signal output
rlabel metal2 s 271694 0 271750 800 6 la_data_out[53]
port 253 nsew signal output
rlabel metal2 s 274730 0 274786 800 6 la_data_out[54]
port 254 nsew signal output
rlabel metal2 s 277766 0 277822 800 6 la_data_out[55]
port 255 nsew signal output
rlabel metal2 s 280802 0 280858 800 6 la_data_out[56]
port 256 nsew signal output
rlabel metal2 s 283838 0 283894 800 6 la_data_out[57]
port 257 nsew signal output
rlabel metal2 s 286874 0 286930 800 6 la_data_out[58]
port 258 nsew signal output
rlabel metal2 s 289910 0 289966 800 6 la_data_out[59]
port 259 nsew signal output
rlabel metal2 s 125966 0 126022 800 6 la_data_out[5]
port 260 nsew signal output
rlabel metal2 s 292946 0 293002 800 6 la_data_out[60]
port 261 nsew signal output
rlabel metal2 s 295982 0 296038 800 6 la_data_out[61]
port 262 nsew signal output
rlabel metal2 s 299018 0 299074 800 6 la_data_out[62]
port 263 nsew signal output
rlabel metal2 s 302054 0 302110 800 6 la_data_out[63]
port 264 nsew signal output
rlabel metal2 s 305090 0 305146 800 6 la_data_out[64]
port 265 nsew signal output
rlabel metal2 s 308126 0 308182 800 6 la_data_out[65]
port 266 nsew signal output
rlabel metal2 s 311162 0 311218 800 6 la_data_out[66]
port 267 nsew signal output
rlabel metal2 s 314198 0 314254 800 6 la_data_out[67]
port 268 nsew signal output
rlabel metal2 s 317234 0 317290 800 6 la_data_out[68]
port 269 nsew signal output
rlabel metal2 s 320270 0 320326 800 6 la_data_out[69]
port 270 nsew signal output
rlabel metal2 s 129002 0 129058 800 6 la_data_out[6]
port 271 nsew signal output
rlabel metal2 s 323306 0 323362 800 6 la_data_out[70]
port 272 nsew signal output
rlabel metal2 s 326342 0 326398 800 6 la_data_out[71]
port 273 nsew signal output
rlabel metal2 s 329378 0 329434 800 6 la_data_out[72]
port 274 nsew signal output
rlabel metal2 s 332414 0 332470 800 6 la_data_out[73]
port 275 nsew signal output
rlabel metal2 s 335450 0 335506 800 6 la_data_out[74]
port 276 nsew signal output
rlabel metal2 s 338486 0 338542 800 6 la_data_out[75]
port 277 nsew signal output
rlabel metal2 s 341522 0 341578 800 6 la_data_out[76]
port 278 nsew signal output
rlabel metal2 s 344558 0 344614 800 6 la_data_out[77]
port 279 nsew signal output
rlabel metal2 s 347594 0 347650 800 6 la_data_out[78]
port 280 nsew signal output
rlabel metal2 s 350630 0 350686 800 6 la_data_out[79]
port 281 nsew signal output
rlabel metal2 s 132038 0 132094 800 6 la_data_out[7]
port 282 nsew signal output
rlabel metal2 s 353666 0 353722 800 6 la_data_out[80]
port 283 nsew signal output
rlabel metal2 s 356702 0 356758 800 6 la_data_out[81]
port 284 nsew signal output
rlabel metal2 s 359738 0 359794 800 6 la_data_out[82]
port 285 nsew signal output
rlabel metal2 s 362774 0 362830 800 6 la_data_out[83]
port 286 nsew signal output
rlabel metal2 s 365810 0 365866 800 6 la_data_out[84]
port 287 nsew signal output
rlabel metal2 s 368846 0 368902 800 6 la_data_out[85]
port 288 nsew signal output
rlabel metal2 s 371882 0 371938 800 6 la_data_out[86]
port 289 nsew signal output
rlabel metal2 s 374918 0 374974 800 6 la_data_out[87]
port 290 nsew signal output
rlabel metal2 s 377954 0 378010 800 6 la_data_out[88]
port 291 nsew signal output
rlabel metal2 s 380990 0 381046 800 6 la_data_out[89]
port 292 nsew signal output
rlabel metal2 s 135074 0 135130 800 6 la_data_out[8]
port 293 nsew signal output
rlabel metal2 s 384026 0 384082 800 6 la_data_out[90]
port 294 nsew signal output
rlabel metal2 s 387062 0 387118 800 6 la_data_out[91]
port 295 nsew signal output
rlabel metal2 s 390098 0 390154 800 6 la_data_out[92]
port 296 nsew signal output
rlabel metal2 s 393134 0 393190 800 6 la_data_out[93]
port 297 nsew signal output
rlabel metal2 s 396170 0 396226 800 6 la_data_out[94]
port 298 nsew signal output
rlabel metal2 s 399206 0 399262 800 6 la_data_out[95]
port 299 nsew signal output
rlabel metal2 s 402242 0 402298 800 6 la_data_out[96]
port 300 nsew signal output
rlabel metal2 s 405278 0 405334 800 6 la_data_out[97]
port 301 nsew signal output
rlabel metal2 s 408314 0 408370 800 6 la_data_out[98]
port 302 nsew signal output
rlabel metal2 s 411350 0 411406 800 6 la_data_out[99]
port 303 nsew signal output
rlabel metal2 s 138110 0 138166 800 6 la_data_out[9]
port 304 nsew signal output
rlabel metal2 s 111798 0 111854 800 6 la_oenb[0]
port 305 nsew signal input
rlabel metal2 s 415398 0 415454 800 6 la_oenb[100]
port 306 nsew signal input
rlabel metal2 s 418434 0 418490 800 6 la_oenb[101]
port 307 nsew signal input
rlabel metal2 s 421470 0 421526 800 6 la_oenb[102]
port 308 nsew signal input
rlabel metal2 s 424506 0 424562 800 6 la_oenb[103]
port 309 nsew signal input
rlabel metal2 s 427542 0 427598 800 6 la_oenb[104]
port 310 nsew signal input
rlabel metal2 s 430578 0 430634 800 6 la_oenb[105]
port 311 nsew signal input
rlabel metal2 s 433614 0 433670 800 6 la_oenb[106]
port 312 nsew signal input
rlabel metal2 s 436650 0 436706 800 6 la_oenb[107]
port 313 nsew signal input
rlabel metal2 s 439686 0 439742 800 6 la_oenb[108]
port 314 nsew signal input
rlabel metal2 s 442722 0 442778 800 6 la_oenb[109]
port 315 nsew signal input
rlabel metal2 s 142158 0 142214 800 6 la_oenb[10]
port 316 nsew signal input
rlabel metal2 s 445758 0 445814 800 6 la_oenb[110]
port 317 nsew signal input
rlabel metal2 s 448794 0 448850 800 6 la_oenb[111]
port 318 nsew signal input
rlabel metal2 s 451830 0 451886 800 6 la_oenb[112]
port 319 nsew signal input
rlabel metal2 s 454866 0 454922 800 6 la_oenb[113]
port 320 nsew signal input
rlabel metal2 s 457902 0 457958 800 6 la_oenb[114]
port 321 nsew signal input
rlabel metal2 s 460938 0 460994 800 6 la_oenb[115]
port 322 nsew signal input
rlabel metal2 s 463974 0 464030 800 6 la_oenb[116]
port 323 nsew signal input
rlabel metal2 s 467010 0 467066 800 6 la_oenb[117]
port 324 nsew signal input
rlabel metal2 s 470046 0 470102 800 6 la_oenb[118]
port 325 nsew signal input
rlabel metal2 s 473082 0 473138 800 6 la_oenb[119]
port 326 nsew signal input
rlabel metal2 s 145194 0 145250 800 6 la_oenb[11]
port 327 nsew signal input
rlabel metal2 s 476118 0 476174 800 6 la_oenb[120]
port 328 nsew signal input
rlabel metal2 s 479154 0 479210 800 6 la_oenb[121]
port 329 nsew signal input
rlabel metal2 s 482190 0 482246 800 6 la_oenb[122]
port 330 nsew signal input
rlabel metal2 s 485226 0 485282 800 6 la_oenb[123]
port 331 nsew signal input
rlabel metal2 s 488262 0 488318 800 6 la_oenb[124]
port 332 nsew signal input
rlabel metal2 s 491298 0 491354 800 6 la_oenb[125]
port 333 nsew signal input
rlabel metal2 s 494334 0 494390 800 6 la_oenb[126]
port 334 nsew signal input
rlabel metal2 s 497370 0 497426 800 6 la_oenb[127]
port 335 nsew signal input
rlabel metal2 s 148230 0 148286 800 6 la_oenb[12]
port 336 nsew signal input
rlabel metal2 s 151266 0 151322 800 6 la_oenb[13]
port 337 nsew signal input
rlabel metal2 s 154302 0 154358 800 6 la_oenb[14]
port 338 nsew signal input
rlabel metal2 s 157338 0 157394 800 6 la_oenb[15]
port 339 nsew signal input
rlabel metal2 s 160374 0 160430 800 6 la_oenb[16]
port 340 nsew signal input
rlabel metal2 s 163410 0 163466 800 6 la_oenb[17]
port 341 nsew signal input
rlabel metal2 s 166446 0 166502 800 6 la_oenb[18]
port 342 nsew signal input
rlabel metal2 s 169482 0 169538 800 6 la_oenb[19]
port 343 nsew signal input
rlabel metal2 s 114834 0 114890 800 6 la_oenb[1]
port 344 nsew signal input
rlabel metal2 s 172518 0 172574 800 6 la_oenb[20]
port 345 nsew signal input
rlabel metal2 s 175554 0 175610 800 6 la_oenb[21]
port 346 nsew signal input
rlabel metal2 s 178590 0 178646 800 6 la_oenb[22]
port 347 nsew signal input
rlabel metal2 s 181626 0 181682 800 6 la_oenb[23]
port 348 nsew signal input
rlabel metal2 s 184662 0 184718 800 6 la_oenb[24]
port 349 nsew signal input
rlabel metal2 s 187698 0 187754 800 6 la_oenb[25]
port 350 nsew signal input
rlabel metal2 s 190734 0 190790 800 6 la_oenb[26]
port 351 nsew signal input
rlabel metal2 s 193770 0 193826 800 6 la_oenb[27]
port 352 nsew signal input
rlabel metal2 s 196806 0 196862 800 6 la_oenb[28]
port 353 nsew signal input
rlabel metal2 s 199842 0 199898 800 6 la_oenb[29]
port 354 nsew signal input
rlabel metal2 s 117870 0 117926 800 6 la_oenb[2]
port 355 nsew signal input
rlabel metal2 s 202878 0 202934 800 6 la_oenb[30]
port 356 nsew signal input
rlabel metal2 s 205914 0 205970 800 6 la_oenb[31]
port 357 nsew signal input
rlabel metal2 s 208950 0 209006 800 6 la_oenb[32]
port 358 nsew signal input
rlabel metal2 s 211986 0 212042 800 6 la_oenb[33]
port 359 nsew signal input
rlabel metal2 s 215022 0 215078 800 6 la_oenb[34]
port 360 nsew signal input
rlabel metal2 s 218058 0 218114 800 6 la_oenb[35]
port 361 nsew signal input
rlabel metal2 s 221094 0 221150 800 6 la_oenb[36]
port 362 nsew signal input
rlabel metal2 s 224130 0 224186 800 6 la_oenb[37]
port 363 nsew signal input
rlabel metal2 s 227166 0 227222 800 6 la_oenb[38]
port 364 nsew signal input
rlabel metal2 s 230202 0 230258 800 6 la_oenb[39]
port 365 nsew signal input
rlabel metal2 s 120906 0 120962 800 6 la_oenb[3]
port 366 nsew signal input
rlabel metal2 s 233238 0 233294 800 6 la_oenb[40]
port 367 nsew signal input
rlabel metal2 s 236274 0 236330 800 6 la_oenb[41]
port 368 nsew signal input
rlabel metal2 s 239310 0 239366 800 6 la_oenb[42]
port 369 nsew signal input
rlabel metal2 s 242346 0 242402 800 6 la_oenb[43]
port 370 nsew signal input
rlabel metal2 s 245382 0 245438 800 6 la_oenb[44]
port 371 nsew signal input
rlabel metal2 s 248418 0 248474 800 6 la_oenb[45]
port 372 nsew signal input
rlabel metal2 s 251454 0 251510 800 6 la_oenb[46]
port 373 nsew signal input
rlabel metal2 s 254490 0 254546 800 6 la_oenb[47]
port 374 nsew signal input
rlabel metal2 s 257526 0 257582 800 6 la_oenb[48]
port 375 nsew signal input
rlabel metal2 s 260562 0 260618 800 6 la_oenb[49]
port 376 nsew signal input
rlabel metal2 s 123942 0 123998 800 6 la_oenb[4]
port 377 nsew signal input
rlabel metal2 s 263598 0 263654 800 6 la_oenb[50]
port 378 nsew signal input
rlabel metal2 s 266634 0 266690 800 6 la_oenb[51]
port 379 nsew signal input
rlabel metal2 s 269670 0 269726 800 6 la_oenb[52]
port 380 nsew signal input
rlabel metal2 s 272706 0 272762 800 6 la_oenb[53]
port 381 nsew signal input
rlabel metal2 s 275742 0 275798 800 6 la_oenb[54]
port 382 nsew signal input
rlabel metal2 s 278778 0 278834 800 6 la_oenb[55]
port 383 nsew signal input
rlabel metal2 s 281814 0 281870 800 6 la_oenb[56]
port 384 nsew signal input
rlabel metal2 s 284850 0 284906 800 6 la_oenb[57]
port 385 nsew signal input
rlabel metal2 s 287886 0 287942 800 6 la_oenb[58]
port 386 nsew signal input
rlabel metal2 s 290922 0 290978 800 6 la_oenb[59]
port 387 nsew signal input
rlabel metal2 s 126978 0 127034 800 6 la_oenb[5]
port 388 nsew signal input
rlabel metal2 s 293958 0 294014 800 6 la_oenb[60]
port 389 nsew signal input
rlabel metal2 s 296994 0 297050 800 6 la_oenb[61]
port 390 nsew signal input
rlabel metal2 s 300030 0 300086 800 6 la_oenb[62]
port 391 nsew signal input
rlabel metal2 s 303066 0 303122 800 6 la_oenb[63]
port 392 nsew signal input
rlabel metal2 s 306102 0 306158 800 6 la_oenb[64]
port 393 nsew signal input
rlabel metal2 s 309138 0 309194 800 6 la_oenb[65]
port 394 nsew signal input
rlabel metal2 s 312174 0 312230 800 6 la_oenb[66]
port 395 nsew signal input
rlabel metal2 s 315210 0 315266 800 6 la_oenb[67]
port 396 nsew signal input
rlabel metal2 s 318246 0 318302 800 6 la_oenb[68]
port 397 nsew signal input
rlabel metal2 s 321282 0 321338 800 6 la_oenb[69]
port 398 nsew signal input
rlabel metal2 s 130014 0 130070 800 6 la_oenb[6]
port 399 nsew signal input
rlabel metal2 s 324318 0 324374 800 6 la_oenb[70]
port 400 nsew signal input
rlabel metal2 s 327354 0 327410 800 6 la_oenb[71]
port 401 nsew signal input
rlabel metal2 s 330390 0 330446 800 6 la_oenb[72]
port 402 nsew signal input
rlabel metal2 s 333426 0 333482 800 6 la_oenb[73]
port 403 nsew signal input
rlabel metal2 s 336462 0 336518 800 6 la_oenb[74]
port 404 nsew signal input
rlabel metal2 s 339498 0 339554 800 6 la_oenb[75]
port 405 nsew signal input
rlabel metal2 s 342534 0 342590 800 6 la_oenb[76]
port 406 nsew signal input
rlabel metal2 s 345570 0 345626 800 6 la_oenb[77]
port 407 nsew signal input
rlabel metal2 s 348606 0 348662 800 6 la_oenb[78]
port 408 nsew signal input
rlabel metal2 s 351642 0 351698 800 6 la_oenb[79]
port 409 nsew signal input
rlabel metal2 s 133050 0 133106 800 6 la_oenb[7]
port 410 nsew signal input
rlabel metal2 s 354678 0 354734 800 6 la_oenb[80]
port 411 nsew signal input
rlabel metal2 s 357714 0 357770 800 6 la_oenb[81]
port 412 nsew signal input
rlabel metal2 s 360750 0 360806 800 6 la_oenb[82]
port 413 nsew signal input
rlabel metal2 s 363786 0 363842 800 6 la_oenb[83]
port 414 nsew signal input
rlabel metal2 s 366822 0 366878 800 6 la_oenb[84]
port 415 nsew signal input
rlabel metal2 s 369858 0 369914 800 6 la_oenb[85]
port 416 nsew signal input
rlabel metal2 s 372894 0 372950 800 6 la_oenb[86]
port 417 nsew signal input
rlabel metal2 s 375930 0 375986 800 6 la_oenb[87]
port 418 nsew signal input
rlabel metal2 s 378966 0 379022 800 6 la_oenb[88]
port 419 nsew signal input
rlabel metal2 s 382002 0 382058 800 6 la_oenb[89]
port 420 nsew signal input
rlabel metal2 s 136086 0 136142 800 6 la_oenb[8]
port 421 nsew signal input
rlabel metal2 s 385038 0 385094 800 6 la_oenb[90]
port 422 nsew signal input
rlabel metal2 s 388074 0 388130 800 6 la_oenb[91]
port 423 nsew signal input
rlabel metal2 s 391110 0 391166 800 6 la_oenb[92]
port 424 nsew signal input
rlabel metal2 s 394146 0 394202 800 6 la_oenb[93]
port 425 nsew signal input
rlabel metal2 s 397182 0 397238 800 6 la_oenb[94]
port 426 nsew signal input
rlabel metal2 s 400218 0 400274 800 6 la_oenb[95]
port 427 nsew signal input
rlabel metal2 s 403254 0 403310 800 6 la_oenb[96]
port 428 nsew signal input
rlabel metal2 s 406290 0 406346 800 6 la_oenb[97]
port 429 nsew signal input
rlabel metal2 s 409326 0 409382 800 6 la_oenb[98]
port 430 nsew signal input
rlabel metal2 s 412362 0 412418 800 6 la_oenb[99]
port 431 nsew signal input
rlabel metal2 s 139122 0 139178 800 6 la_oenb[9]
port 432 nsew signal input
rlabel metal4 s 4208 2128 4528 297616 6 vccd1
port 433 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 297616 6 vccd1
port 433 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 297616 6 vccd1
port 433 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 297616 6 vccd1
port 433 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 297616 6 vccd1
port 433 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 297616 6 vccd1
port 433 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 297616 6 vccd1
port 433 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 297616 6 vccd1
port 433 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 297616 6 vccd1
port 433 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 297616 6 vccd1
port 433 nsew power bidirectional
rlabel metal4 s 311408 2128 311728 297616 6 vccd1
port 433 nsew power bidirectional
rlabel metal4 s 342128 2128 342448 297616 6 vccd1
port 433 nsew power bidirectional
rlabel metal4 s 372848 2128 373168 297616 6 vccd1
port 433 nsew power bidirectional
rlabel metal4 s 403568 2128 403888 297616 6 vccd1
port 433 nsew power bidirectional
rlabel metal4 s 434288 2128 434608 297616 6 vccd1
port 433 nsew power bidirectional
rlabel metal4 s 465008 2128 465328 297616 6 vccd1
port 433 nsew power bidirectional
rlabel metal4 s 495728 2128 496048 297616 6 vccd1
port 433 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 297616 6 vssd1
port 434 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 297616 6 vssd1
port 434 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 297616 6 vssd1
port 434 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 297616 6 vssd1
port 434 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 297616 6 vssd1
port 434 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 297616 6 vssd1
port 434 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 297616 6 vssd1
port 434 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 297616 6 vssd1
port 434 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 297616 6 vssd1
port 434 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 297616 6 vssd1
port 434 nsew ground bidirectional
rlabel metal4 s 326768 2128 327088 297616 6 vssd1
port 434 nsew ground bidirectional
rlabel metal4 s 357488 2128 357808 297616 6 vssd1
port 434 nsew ground bidirectional
rlabel metal4 s 388208 2128 388528 297616 6 vssd1
port 434 nsew ground bidirectional
rlabel metal4 s 418928 2128 419248 297616 6 vssd1
port 434 nsew ground bidirectional
rlabel metal4 s 449648 2128 449968 297616 6 vssd1
port 434 nsew ground bidirectional
rlabel metal4 s 480368 2128 480688 297616 6 vssd1
port 434 nsew ground bidirectional
rlabel metal2 s 2502 0 2558 800 6 wb_ack
port 435 nsew signal output
rlabel metal2 s 8574 0 8630 800 6 wb_addr_i[0]
port 436 nsew signal input
rlabel metal2 s 38934 0 38990 800 6 wb_addr_i[10]
port 437 nsew signal input
rlabel metal2 s 41970 0 42026 800 6 wb_addr_i[11]
port 438 nsew signal input
rlabel metal2 s 45006 0 45062 800 6 wb_addr_i[12]
port 439 nsew signal input
rlabel metal2 s 48042 0 48098 800 6 wb_addr_i[13]
port 440 nsew signal input
rlabel metal2 s 51078 0 51134 800 6 wb_addr_i[14]
port 441 nsew signal input
rlabel metal2 s 54114 0 54170 800 6 wb_addr_i[15]
port 442 nsew signal input
rlabel metal2 s 57150 0 57206 800 6 wb_addr_i[16]
port 443 nsew signal input
rlabel metal2 s 60186 0 60242 800 6 wb_addr_i[17]
port 444 nsew signal input
rlabel metal2 s 63222 0 63278 800 6 wb_addr_i[18]
port 445 nsew signal input
rlabel metal2 s 66258 0 66314 800 6 wb_addr_i[19]
port 446 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 wb_addr_i[1]
port 447 nsew signal input
rlabel metal2 s 69294 0 69350 800 6 wb_addr_i[20]
port 448 nsew signal input
rlabel metal2 s 72330 0 72386 800 6 wb_addr_i[21]
port 449 nsew signal input
rlabel metal2 s 75366 0 75422 800 6 wb_addr_i[22]
port 450 nsew signal input
rlabel metal2 s 78402 0 78458 800 6 wb_addr_i[23]
port 451 nsew signal input
rlabel metal2 s 81438 0 81494 800 6 wb_addr_i[24]
port 452 nsew signal input
rlabel metal2 s 84474 0 84530 800 6 wb_addr_i[25]
port 453 nsew signal input
rlabel metal2 s 87510 0 87566 800 6 wb_addr_i[26]
port 454 nsew signal input
rlabel metal2 s 90546 0 90602 800 6 wb_addr_i[27]
port 455 nsew signal input
rlabel metal2 s 93582 0 93638 800 6 wb_addr_i[28]
port 456 nsew signal input
rlabel metal2 s 96618 0 96674 800 6 wb_addr_i[29]
port 457 nsew signal input
rlabel metal2 s 14646 0 14702 800 6 wb_addr_i[2]
port 458 nsew signal input
rlabel metal2 s 99654 0 99710 800 6 wb_addr_i[30]
port 459 nsew signal input
rlabel metal2 s 102690 0 102746 800 6 wb_addr_i[31]
port 460 nsew signal input
rlabel metal2 s 17682 0 17738 800 6 wb_addr_i[3]
port 461 nsew signal input
rlabel metal2 s 20718 0 20774 800 6 wb_addr_i[4]
port 462 nsew signal input
rlabel metal2 s 23754 0 23810 800 6 wb_addr_i[5]
port 463 nsew signal input
rlabel metal2 s 26790 0 26846 800 6 wb_addr_i[6]
port 464 nsew signal input
rlabel metal2 s 29826 0 29882 800 6 wb_addr_i[7]
port 465 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 wb_addr_i[8]
port 466 nsew signal input
rlabel metal2 s 35898 0 35954 800 6 wb_addr_i[9]
port 467 nsew signal input
rlabel metal2 s 3514 0 3570 800 6 wb_clk_i
port 468 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 wb_cyc_i
port 469 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 wb_data_i[0]
port 470 nsew signal input
rlabel metal2 s 39946 0 40002 800 6 wb_data_i[10]
port 471 nsew signal input
rlabel metal2 s 42982 0 43038 800 6 wb_data_i[11]
port 472 nsew signal input
rlabel metal2 s 46018 0 46074 800 6 wb_data_i[12]
port 473 nsew signal input
rlabel metal2 s 49054 0 49110 800 6 wb_data_i[13]
port 474 nsew signal input
rlabel metal2 s 52090 0 52146 800 6 wb_data_i[14]
port 475 nsew signal input
rlabel metal2 s 55126 0 55182 800 6 wb_data_i[15]
port 476 nsew signal input
rlabel metal2 s 58162 0 58218 800 6 wb_data_i[16]
port 477 nsew signal input
rlabel metal2 s 61198 0 61254 800 6 wb_data_i[17]
port 478 nsew signal input
rlabel metal2 s 64234 0 64290 800 6 wb_data_i[18]
port 479 nsew signal input
rlabel metal2 s 67270 0 67326 800 6 wb_data_i[19]
port 480 nsew signal input
rlabel metal2 s 12622 0 12678 800 6 wb_data_i[1]
port 481 nsew signal input
rlabel metal2 s 70306 0 70362 800 6 wb_data_i[20]
port 482 nsew signal input
rlabel metal2 s 73342 0 73398 800 6 wb_data_i[21]
port 483 nsew signal input
rlabel metal2 s 76378 0 76434 800 6 wb_data_i[22]
port 484 nsew signal input
rlabel metal2 s 79414 0 79470 800 6 wb_data_i[23]
port 485 nsew signal input
rlabel metal2 s 82450 0 82506 800 6 wb_data_i[24]
port 486 nsew signal input
rlabel metal2 s 85486 0 85542 800 6 wb_data_i[25]
port 487 nsew signal input
rlabel metal2 s 88522 0 88578 800 6 wb_data_i[26]
port 488 nsew signal input
rlabel metal2 s 91558 0 91614 800 6 wb_data_i[27]
port 489 nsew signal input
rlabel metal2 s 94594 0 94650 800 6 wb_data_i[28]
port 490 nsew signal input
rlabel metal2 s 97630 0 97686 800 6 wb_data_i[29]
port 491 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 wb_data_i[2]
port 492 nsew signal input
rlabel metal2 s 100666 0 100722 800 6 wb_data_i[30]
port 493 nsew signal input
rlabel metal2 s 103702 0 103758 800 6 wb_data_i[31]
port 494 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 wb_data_i[3]
port 495 nsew signal input
rlabel metal2 s 21730 0 21786 800 6 wb_data_i[4]
port 496 nsew signal input
rlabel metal2 s 24766 0 24822 800 6 wb_data_i[5]
port 497 nsew signal input
rlabel metal2 s 27802 0 27858 800 6 wb_data_i[6]
port 498 nsew signal input
rlabel metal2 s 30838 0 30894 800 6 wb_data_i[7]
port 499 nsew signal input
rlabel metal2 s 33874 0 33930 800 6 wb_data_i[8]
port 500 nsew signal input
rlabel metal2 s 36910 0 36966 800 6 wb_data_i[9]
port 501 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 wb_data_o[0]
port 502 nsew signal output
rlabel metal2 s 40958 0 41014 800 6 wb_data_o[10]
port 503 nsew signal output
rlabel metal2 s 43994 0 44050 800 6 wb_data_o[11]
port 504 nsew signal output
rlabel metal2 s 47030 0 47086 800 6 wb_data_o[12]
port 505 nsew signal output
rlabel metal2 s 50066 0 50122 800 6 wb_data_o[13]
port 506 nsew signal output
rlabel metal2 s 53102 0 53158 800 6 wb_data_o[14]
port 507 nsew signal output
rlabel metal2 s 56138 0 56194 800 6 wb_data_o[15]
port 508 nsew signal output
rlabel metal2 s 59174 0 59230 800 6 wb_data_o[16]
port 509 nsew signal output
rlabel metal2 s 62210 0 62266 800 6 wb_data_o[17]
port 510 nsew signal output
rlabel metal2 s 65246 0 65302 800 6 wb_data_o[18]
port 511 nsew signal output
rlabel metal2 s 68282 0 68338 800 6 wb_data_o[19]
port 512 nsew signal output
rlabel metal2 s 13634 0 13690 800 6 wb_data_o[1]
port 513 nsew signal output
rlabel metal2 s 71318 0 71374 800 6 wb_data_o[20]
port 514 nsew signal output
rlabel metal2 s 74354 0 74410 800 6 wb_data_o[21]
port 515 nsew signal output
rlabel metal2 s 77390 0 77446 800 6 wb_data_o[22]
port 516 nsew signal output
rlabel metal2 s 80426 0 80482 800 6 wb_data_o[23]
port 517 nsew signal output
rlabel metal2 s 83462 0 83518 800 6 wb_data_o[24]
port 518 nsew signal output
rlabel metal2 s 86498 0 86554 800 6 wb_data_o[25]
port 519 nsew signal output
rlabel metal2 s 89534 0 89590 800 6 wb_data_o[26]
port 520 nsew signal output
rlabel metal2 s 92570 0 92626 800 6 wb_data_o[27]
port 521 nsew signal output
rlabel metal2 s 95606 0 95662 800 6 wb_data_o[28]
port 522 nsew signal output
rlabel metal2 s 98642 0 98698 800 6 wb_data_o[29]
port 523 nsew signal output
rlabel metal2 s 16670 0 16726 800 6 wb_data_o[2]
port 524 nsew signal output
rlabel metal2 s 101678 0 101734 800 6 wb_data_o[30]
port 525 nsew signal output
rlabel metal2 s 104714 0 104770 800 6 wb_data_o[31]
port 526 nsew signal output
rlabel metal2 s 19706 0 19762 800 6 wb_data_o[3]
port 527 nsew signal output
rlabel metal2 s 22742 0 22798 800 6 wb_data_o[4]
port 528 nsew signal output
rlabel metal2 s 25778 0 25834 800 6 wb_data_o[5]
port 529 nsew signal output
rlabel metal2 s 28814 0 28870 800 6 wb_data_o[6]
port 530 nsew signal output
rlabel metal2 s 31850 0 31906 800 6 wb_data_o[7]
port 531 nsew signal output
rlabel metal2 s 34886 0 34942 800 6 wb_data_o[8]
port 532 nsew signal output
rlabel metal2 s 37922 0 37978 800 6 wb_data_o[9]
port 533 nsew signal output
rlabel metal2 s 5538 0 5594 800 6 wb_rst_i
port 534 nsew signal input
rlabel metal2 s 6550 0 6606 800 6 wb_stb
port 535 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 wb_we_i
port 536 nsew signal input
rlabel metal2 s 105726 0 105782 800 6 wbs_sel_i[0]
port 537 nsew signal input
rlabel metal2 s 106738 0 106794 800 6 wbs_sel_i[1]
port 538 nsew signal input
rlabel metal2 s 107750 0 107806 800 6 wbs_sel_i[2]
port 539 nsew signal input
rlabel metal2 s 108762 0 108818 800 6 wbs_sel_i[3]
port 540 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 500000 300000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 38979316
string GDS_FILE /home/leviathan/kicp/openlane/AI_Accelerator_Top/runs/23_06_03_19_49/results/signoff/AI_Accelerator_Top.magic.gds
string GDS_START 220712
<< end >>

